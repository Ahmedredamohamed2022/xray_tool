** NOTE: ngspice DOES NOT handle environment variables used in the test benches. the Makefile handles that for you, if you wish to use your own command make sure you manually update the spice files
VSS2 VSS GND 0
.save i(VSS2)
vtot net1 VDD 0
.save i(vtot)
VDD1 EN VSS 1.8
.save i(VDD1)
VDD2 net1 VSS ${VDD_VAL}
.save i(VDD2)


x1 VOUT VIP EN VOUT VDD VSS EF_AMP3V3
 
VDD4 VIP VSS sin(1.65 ${VPEAK} ${FREQ})
.save i(VDD4)
C1 VOUT VSS 5p m=1
R1 VOUT net2 10k m=1

.options RSHUNT=1e15
.options savecurrents
.option TEMP=${TEMP_VAL}
.option TNOM=${TEMP_VAL}
.option interp
.control
set wr_singlescale
set wr_vecnames
declare thd_VOUT
**set filetype=binary
set filetype=ascii
set color0=white
set color1=black
set color3=blue
set xbrushwidth=3
save all
run
op
tran ${T_START} ${T_STOP} ${T_STEP}
*tran 0.001u 0.002m 0.010u
let vi=v(VIP)-1.65
let VOUT=v(VOUT)-1.65
 

fourier ${FREQ} vi VOUT
let idx = 2
let sum_mag_square = 0
while idx < 10
    let mag = fourier11[1][idx]
    let sum_mag_square = sum_mag_square + mag * mag
    let idx = idx + 1
end
let root_sum_mag_square = sqrt(sum_mag_square)
let thd_vi = root_sum_mag_square / fourier11[1][1] * 100
print thd_vi

let idx = 2
let sum_mag_square = 0
while idx < 10
    let mag = fourier12[1][idx]
    let sum_mag_square = sum_mag_square + mag * mag
    let idx = idx + 1
end
let root_sum_mag_square = sqrt(sum_mag_square)
let thd_VOUT = root_sum_mag_square / fourier12[1][1] * 100
print thd_VOUT


let pvt_c=${ENUMER_CASE_NBR}+1
let VDD_VAL=${VDD_VAL} 
let DVDD_VAL=${DVDD_VAL} 
let TEMP_VAL=${TEMP_VAL}

echo "TEMP ${TEMP_VAL} VDD ${VDD_VAL} DVDD ${DVDD_VAL} e:${ENUMER_CASE_NBR}_tran:${CORNERS}_temp:${TEMP_VAL}_VDD:${VDD_VAL}" "thd_VOUT" $&thd_VOUT  eol  >> out.txt	   
write /ciic/designs/analog-mixed-signal-blocks/Xschem-schematic/EF_AMP3V3/xray/ampthdpvt/rawfiles-enumer/e:${ENUMER_CASE_NBR}_temp:${TEMP_VAL}__VDD:${VDD_VAL}_DVDD:${DVDD_VAL}_tran:${CORNERS}.raw 
+ {thd_VOUT}  {VDD_VAL}  {DVDD_VAL}  {TEMP_VAL}
write /ciic/designs/analog-mixed-signal-blocks/Xschem-schematic/EF_AMP3V3/xray/ampthdpvt/rawfiles/pvt{$&pvt_c}.raw 
+ {thd_VOUT}  {VDD_VAL}  {DVDD_VAL}  {TEMP_VAL}

.endc


.include /ciic/pdk//sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice
.include /ciic/pdk//sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice
.lib /ciic/pdk//sky130A/libs.tech/ngspice/sky130.lib.spice ${CORNERS}
.include /ciic/designs/analog-mixed-signal-blocks/Xschem-schematic/EF_AMP3V3/xray/EF_AMP3V3.spice




.GLOBAL GND
.end
