** sch_path:
*+ /ciic/designs/analog-mixed-signal-blocks/Xschem-schematic/ota-2stage/ndiff-ota/tb-ac-openloop/openloopgain-psneg.sch
**.subckt openloopgain-psneg
V1 vss GND 0 ac=1
V2 vdd vss ${VDD} ac=0
I0 vdd ibiasn ${IBIASN}
V3 vip net1 ${VCOM}
V4 vin net1 ${VCOM}
X1 vout vdd vss ibiasn vip vin ndiff-ota-circuit
V5 net1 vss 0 ac=0
C1 vout vss ${CL} m=1
**** begin user architecture code
.lib /ciic/pdk//sky130A/libs.tech/ngspice/sky130.lib.spice ${CORNERS}
.control
**set filetype=binary
set filetype=ascii
ac dec ${ND} ${FSTART} ${FSTOP}
set units = degrees
set color0=white
set color1=black
set color3=blue
set xbrushwidth=3
plot db(vout) phase(vout)
meas ac psnegr FIND vdb(vout) AT=10
echo  $&psnegr  >> psneg.txt
write  /ciic/designs/analog-mixed-signal-blocks/Xschem-schematic/ota-2stage/xray4ota/ac/psneg/rawfiles/psneggain.raw
+   {psnegr}
.endc
.end
.GLOBAL GND
.end
