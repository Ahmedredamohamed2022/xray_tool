* NGSPICE file created from EF_AMP3V3.ext - technology: sky130A

.subckt EF_AMP3V3 VOUT VIP EN VIN VDD VSS
X0 VOUT.t338 pdrv1.t2 VDD.t368 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X1 VOUT.t337 pdrv1.t3 VDD.t367 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X2 VOUT.t38 ndrv.t0 VSS.t137 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X3 VOUT.t336 pdrv1.t4 VDD.t366 VDD.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X4 VDD.t370 pdrv2.t0 VOUT.t342 VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X5 VOUT.t335 pdrv1.t5 VDD.t365 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X6 VDD.t152 pdrv2.t1 VOUT.t126 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X7 VDD.t153 pdrv2.t2 VOUT.t127 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X8 VDD.t162 a_n1922_640# pdrv1.t1 VDD.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X9 VOUT.t334 pdrv1.t6 VDD.t364 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X10 VDD.t363 pdrv1.t7 VOUT.t333 VDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X11 VSS.t136 ndrv.t1 VOUT.t382 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X12 VOUT.t88 pdrv2.t3 VDD.t109 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X13 VOUT.t332 pdrv1.t8 VDD.t362 VDD.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X14 VOUT.t418 pdrv2.t4 VDD.t419 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X15 VDD.t108 pdrv2.t5 VOUT.t87 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X16 VDD.t414 pdrv2.t6 VOUT.t406 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X17 VOUT.t472 ndrv.t2 VSS.t135 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X18 VOUT.t478 pdrv2.t7 VDD.t436 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X19 VDD.t361 pdrv1.t9 VOUT.t331 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X20 VOUT.t17 pdrv2.t8 VDD.t14 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X21 VOUT.t464 pdrv2.t9 VDD.t434 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X22 VDD.t360 pdrv1.t10 VOUT.t330 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X23 VSS.t134 ndrv.t3 VOUT.t467 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X24 VOUT.t329 pdrv1.t11 VDD.t359 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X25 VDD.t151 pdrv2.t10 VOUT.t125 VDD.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X26 VOUT.t328 pdrv1.t12 VDD.t358 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X27 VSS.t133 ndrv.t4 VOUT.t476 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X28 nbias.t7 nbias.t6 VSS.t9 VSS.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X29 VDD.t46 pdrv2.t11 VOUT.t37 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X30 VOUT.t397 pdrv2.t12 VDD.t411 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X31 VOUT.t327 pdrv1.t13 VDD.t357 VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X32 VDD.t376 pdrv2.t13 VOUT.t352 VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X33 VOUT.t326 pdrv1.t14 VDD.t356 VDD.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X34 VOUT.t2 ndrv.t5 VSS.t132 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X35 VDD.t355 pdrv1.t15 VOUT.t325 VDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X36 VDD.t354 pdrv1.t16 VOUT.t324 VDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X37 VOUT.t383 ndrv.t6 VSS.t131 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X38 VDD.t410 pdrv2.t14 VOUT.t395 VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X39 VOUT.t97 ndrv.t7 VSS.t130 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X40 VOUT.t323 pdrv1.t17 VDD.t353 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X41 VDD.t154 pdrv2.t15 VOUT.t129 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X42 VOUT.t322 pdrv1.t18 VDD.t352 VDD.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X43 VDD.t429 pdrv2.t16 VOUT.t438 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X44 VDD.t409 pdrv2.t17 VOUT.t394 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X45 VOUT.t18 pdrv2.t18 VDD.t16 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X46 VDD.t351 pdrv1.t19 VOUT.t321 VDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X47 VDD.t350 pdrv1.t20 VOUT.t320 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X48 VOUT.t319 pdrv1.t21 VDD.t349 VDD.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X49 VOUT.t340 pdrv2.t19 VDD.t369 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X50 VOUT.t350 pdrv2.t20 VDD.t374 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X51 VDD.t448 pdrv2.t21 VOUT.t494 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X52 VOUT.t109 pdrv2.t22 VDD.t132 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X53 VOUT.t413 pdrv2.t23 VDD.t416 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X54 VOUT.t318 pdrv1.t22 VDD.t344 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X55 VSS.t129 ndrv.t8 VOUT.t339 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X56 VDD.t348 pdrv1.t23 VOUT.t317 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X57 VOUT.t316 pdrv1.t24 VDD.t347 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X58 VDD.t346 pdrv1.t25 VOUT.t315 VDD.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X59 VSS.t128 ndrv.t9 VOUT.t469 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X60 VOUT.t314 pdrv1.t26 VDD.t345 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X61 VOUT.t29 pdrv2.t24 VDD.t41 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X62 VDD.t343 pdrv1.t27 VOUT.t313 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X63 VDD.t397 pdrv2.t25 VOUT.t377 VDD.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X64 VOUT.t312 pdrv1.t28 VDD.t342 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X65 VDD.t426 pdrv2.t26 VOUT.t428 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X66 VSS.t127 ndrv.t10 VOUT.t456 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X67 VOUT.t311 pdrv1.t29 VDD.t341 VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X68 VOUT.t310 pdrv1.t30 VDD.t340 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X69 VOUT.t415 pdrv2.t27 VDD.t418 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X70 VSS.t126 ndrv.t11 VOUT.t455 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X71 VOUT.t309 pdrv1.t31 VDD.t339 VDD.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X72 VDD.t423 pdrv2.t28 VOUT.t423 VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X73 VOUT.t461 ndrv.t12 VSS.t125 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X74 VOUT.t42 pdrv2.t29 VDD.t52 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X75 VDD.t338 pdrv1.t32 VOUT.t308 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X76 VDD.t337 pdrv1.t33 VOUT.t307 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X77 a_n3090_640# VIN.t0 vcomn2 VSS.t1 sky130_fd_pr__nfet_03v3_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X78 VSS.t124 ndrv.t13 VOUT.t468 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X79 VDD.t420 pdrv2.t30 VOUT.t419 VDD.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X80 VOUT.t306 pdrv1.t34 VDD.t336 VDD.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X81 VDD.t335 pdrv1.t35 VOUT.t305 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X82 VDD.t334 pdrv1.t36 VOUT.t304 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X83 pdrv1.t1 a_n1922_640# VDD.t160 VDD.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X84 VOUT.t12 pdrv2.t31 VDD.t10 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X85 a_n1922_640# VIN.t1 vcomn1 VSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X86 VDD.t40 pbias vcomp VDD.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X87 VDD.t333 pdrv1.t37 VOUT.t303 VDD.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X88 VSS.t123 ndrv.t14 VOUT.t477 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X89 VOUT.t302 pdrv1.t38 VDD.t332 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X90 VOUT.t301 pdrv1.t39 VDD.t331 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X91 VOUT.t300 pdrv1.t40 VDD.t330 VDD.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X92 VOUT.t299 pdrv1.t41 VDD.t329 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X93 VSS.t122 ndrv.t15 VOUT.t480 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X94 VOUT.t298 pdrv1.t42 VDD.t328 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X95 VDD.t327 pdrv1.t43 VOUT.t297 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X96 VDD.t407 pdrv2.t32 VOUT.t391 VDD.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X97 VOUT.t296 pdrv1.t44 VDD.t326 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X98 VSS.t121 ndrv.t16 VOUT.t475 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X99 VOUT.t295 pdrv1.t45 VDD.t325 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X100 VDD.t324 pdrv1.t46 VOUT.t294 VDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X101 VDD.t421 pdrv2.t33 VOUT.t421 VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X102 VSS.t120 ndrv.t17 VOUT.t457 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X103 VOUT.t293 pdrv1.t47 VDD.t323 VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X104 VOUT.t1 ndrv.t18 VSS.t119 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X105 VOUT.t292 pdrv1.t48 VDD.t322 VDD.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X106 VSS.t118 ndrv.t19 VOUT.t448 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X107 VDD.t321 pdrv1.t49 VOUT.t291 VDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X108 VDD.t12 pdrv2.t34 VOUT.t13 VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X109 VOUT.t454 ndrv.t20 VSS.t117 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X110 VDD.t417 pdrv2.t35 VOUT.t414 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X111 VOUT.t401 ndrv.t21 VSS.t116 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X112 VDD.t111 pdrv2.t36 VOUT.t90 VDD.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X113 VOUT.t460 ndrv.t22 VSS.t115 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X114 VOUT.t483 pdrv2.t37 VDD.t437 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X115 a_n551_n345# VIN.t2 vcomp VDD.t446 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X116 VOUT.t290 pdrv1.t50 VDD.t320 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X117 VSS.t114 ndrv.t23 VOUT.t459 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X118 VDD.t319 pdrv1.t51 VOUT.t289 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X119 VOUT.t288 pdrv1.t52 VDD.t318 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X120 VDD.t317 pdrv1.t53 VOUT.t287 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X121 VOUT.t458 ndrv.t24 VSS.t113 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X122 VOUT.t427 pdrv2.t38 VDD.t425 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X123 VOUT.t449 ndrv.t25 VSS.t112 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X124 VSS.t111 ndrv.t26 VOUT.t403 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X125 VOUT.t484 ndrv.t27 VSS.t110 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X126 VOUT.t381 pdrv2.t39 VDD.t400 VDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X127 VOUT.t447 ndrv.t28 VSS.t109 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X128 VOUT.t466 pdrv2.t40 VDD.t435 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X129 vcomp pbias VDD.t38 VDD.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X130 VDD.t316 pdrv1.t54 VOUT.t286 VDD.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X131 VOUT.t285 pdrv1.t55 VDD.t315 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X132 VDD.t427 pdrv2.t41 VOUT.t429 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X133 VSS.t108 ndrv.t29 VOUT.t453 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X134 VOUT.t284 pdrv1.t56 VDD.t314 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X135 VOUT.t452 ndrv.t30 VSS.t107 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X136 VDD.t313 pdrv1.t57 VOUT.t283 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X137 VSS.t106 ndrv.t31 VOUT.t451 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X138 VDD.t87 pdrv2.t42 VOUT.t70 VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X139 VDD.t415 pdrv2.t43 VOUT.t412 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X140 VSS.t105 ndrv.t32 VOUT.t450 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X141 VOUT.t282 pdrv1.t58 VDD.t312 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X142 VDD.t131 pdrv2.t44 VOUT.t107 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X143 VOUT.t482 ndrv.t33 VSS.t104 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X144 VDD.t311 pdrv1.t59 VOUT.t281 VDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X145 VOUT.t135 ndrv.t34 VSS.t103 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X146 VOUT.t280 pdrv1.t60 VDD.t310 VDD.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X147 VOUT.t425 pdrv2.t45 VDD.t424 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X148 VDD.t306 pdrv1.t61 VOUT.t279 VDD.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X149 VOUT.t433 ndrv.t35 VSS.t102 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X150 VOUT.t518 ndrv.t36 VSS.t101 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X151 VSS.t100 ndrv.t37 VOUT.t446 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X152 VDD.t309 pdrv1.t62 VOUT.t278 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X153 VOUT.t363 pdrv2.t46 VDD.t383 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X154 VDD.t308 pdrv1.t63 VOUT.t277 VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X155 VOUT.t445 ndrv.t38 VSS.t99 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X156 VDD.t412 pdrv2.t47 VOUT.t404 VDD.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X157 VDD.t307 pdrv1.t64 VOUT.t276 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X158 VDD.t305 pdrv1.t65 VOUT.t275 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X159 VDD.t125 pdrv2.t48 VOUT.t102 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X160 VOUT.t274 pdrv1.t66 VDD.t304 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X161 VOUT.t273 pdrv1.t67 VDD.t303 VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X162 VOUT.t272 pdrv1.t68 VDD.t302 VDD.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X163 VOUT.t51 pdrv2.t49 VDD.t67 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X164 VSS.t98 ndrv.t39 VOUT.t444 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X165 VDD.t9 pdrv2.t50 VOUT.t9 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X166 VSS.t97 ndrv.t40 VOUT.t443 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X167 VOUT.t271 pdrv1.t69 VDD.t297 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X168 VDD.t301 pdrv1.t70 VOUT.t270 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X169 VOUT.t269 pdrv1.t71 VDD.t300 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X170 VDD.t299 pdrv1.t72 VOUT.t268 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X171 VOUT.t267 pdrv1.t73 VDD.t298 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X172 VOUT.t266 pdrv1.t74 VDD.t296 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X173 VOUT.t265 pdrv1.t75 VDD.t295 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X174 VSS.t96 ndrv.t41 VOUT.t434 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X175 VDD.t127 pdrv2.t51 VOUT.t104 VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X176 VDD.t294 pdrv1.t76 VOUT.t264 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X177 VDD.t466 pdrv2.t52 VOUT.t513 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X178 VDD.t106 pdrv2.t53 VOUT.t85 VDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X179 VOUT.t137 ndrv.t42 VSS.t95 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X180 VOUT.t138 ndrv.t43 VSS.t94 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X181 VDD.t293 pdrv1.t77 VOUT.t263 VDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X182 VSS.t93 ndrv.t44 VOUT.t10 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X183 VDD.t292 pdrv1.t78 VOUT.t262 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X184 VDD.t431 pdrv2.t54 VOUT.t441 VDD.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X185 VOUT.t261 pdrv1.t79 VDD.t291 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X186 VDD.t413 pdrv2.t55 VOUT.t405 VDD.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X187 VSS.t92 ndrv.t45 VOUT.t515 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X188 VSS.t91 ndrv.t46 VOUT.t514 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X189 VOUT.t19 pdrv2.t56 VDD.t18 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X190 VOUT.t11 ndrv.t47 VSS.t90 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X191 VDD.t290 pdrv1.t80 VOUT.t260 VDD.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X192 VOUT.t136 ndrv.t48 VSS.t89 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X193 VDD.t289 pdrv1.t81 VOUT.t259 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X194 VOUT.t258 pdrv1.t82 VDD.t288 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X195 VDD.t287 pdrv1.t83 VOUT.t257 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X196 VOUT.t50 ndrv.t49 VSS.t88 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X197 VOUT.t34 pdrv2.t57 VDD.t44 VDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X198 VOUT.t56 pdrv2.t58 VDD.t69 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X199 VOUT.t35 ndrv.t50 VSS.t87 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X200 nbias.t5 nbias.t4 VSS.t6 VSS.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X201 VOUT.t256 pdrv1.t84 VDD.t286 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X202 VDD.t285 pdrv1.t85 VOUT.t255 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X203 VDD.t95 pdrv2.t59 VOUT.t75 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X204 VDD.t68 pdrv2.t60 VOUT.t52 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X205 VOUT.t254 pdrv1.t86 VDD.t284 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X206 VOUT.t485 pdrv2.t61 VDD.t438 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X207 VDD.t283 pdrv1.t87 VOUT.t253 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X208 VOUT.t252 pdrv1.t88 VDD.t282 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X209 VDD.t126 pdrv2.t62 VOUT.t103 VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X210 VOUT.t251 pdrv1.t89 VDD.t281 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X211 VDD.t130 pdrv2.t63 VOUT.t106 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X212 VOUT.t402 ndrv.t51 VSS.t86 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X213 VOUT.t250 pdrv1.t90 VDD.t280 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X214 VDD.t371 pdrv2.t64 VOUT.t343 VDD.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X215 VOUT.t60 ndrv.t52 VSS.t85 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X216 VOUT.t440 pdrv2.t65 VDD.t430 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X217 VDD.t279 pdrv1.t91 VOUT.t249 VDD.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X218 VSS.t84 ndrv.t53 VOUT.t0 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X219 VOUT.t248 pdrv1.t92 VDD.t278 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X220 VDD.t277 pdrv1.t93 VOUT.t247 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X221 VDD.t276 pdrv1.t94 VOUT.t246 VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X222 VOUT.t349 pdrv2.t66 VDD.t373 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X223 VDD.t408 pdrv2.t67 VOUT.t393 VDD.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X224 VSS.t83 ndrv.t54 VOUT.t435 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X225 VOUT.t32 pdrv2.t68 VDD.t43 VDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X226 VOUT.t436 ndrv.t55 VSS.t82 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X227 VDD.t158 a_n1922_640# a_n1922_640# VDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X228 VOUT.t245 pdrv1.t95 VDD.t275 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X229 VDD.t274 pdrv1.t96 VOUT.t244 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X230 VDD.t273 pdrv1.t97 VOUT.t243 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X231 VDD.t422 pdrv2.t69 VOUT.t422 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X232 a_n551_n345# a_n551_n345# VSS.t4 VSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X233 VOUT.t242 pdrv1.t98 VDD.t272 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X234 VSS.t81 ndrv.t56 VOUT.t84 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X235 VDD.t107 pdrv2.t70 VOUT.t86 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X236 VDD.t271 pdrv1.t99 VOUT.t241 VDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X237 VOUT.t101 pdrv2.t71 VDD.t124 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X238 VSS.t80 ndrv.t57 VOUT.t16 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X239 VOUT.t41 pdrv2.t72 VDD.t51 VDD.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X240 VDD.t112 pdrv2.t73 VOUT.t91 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X241 VOUT.t240 pdrv1.t100 VDD.t270 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X242 VDD.t269 pdrv1.t101 VOUT.t239 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X243 VOUT.t238 pdrv1.t102 VDD.t268 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X244 VDD.t433 pdrv2.t74 VOUT.t463 VDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X245 VOUT.t237 pdrv1.t103 VDD.t267 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X246 VOUT.t8 pdrv2.t75 VDD.t7 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X247 VOUT.t398 ndrv.t58 VSS.t79 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X248 VDD.t375 pdrv2.t76 VOUT.t351 VDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X249 VDD.t266 pdrv1.t104 VOUT.t236 VDD.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X250 VDD.t428 pdrv2.t77 VOUT.t430 VDD.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X251 VSS.t78 ndrv.t59 VOUT.t108 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X252 VOUT.t235 pdrv1.t105 VDD.t265 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X253 VDD.t264 pdrv1.t106 VOUT.t234 VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X254 VDD.t263 pdrv1.t107 VOUT.t233 VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X255 VOUT.t353 pdrv2.t78 VDD.t377 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X256 VDD.t432 pdrv2.t79 VOUT.t462 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X257 VDD.t262 pdrv1.t108 VOUT.t232 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X258 VDD.t388 pdrv2.t80 VOUT.t368 VDD.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X259 VDD.t381 pdrv2.t81 VOUT.t358 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X260 VOUT.t132 pdrv2.t82 VDD.t165 VDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X261 VOUT.t437 ndrv.t60 VSS.t77 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X262 VDD.t261 pdrv1.t109 VOUT.t231 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X263 VOUT.t399 ndrv.t61 VSS.t76 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X264 VOUT.t230 pdrv1.t110 VDD.t260 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X265 VOUT.t229 pdrv1.t111 VDD.t259 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X266 VOUT.t27 pdrv2.t83 VDD.t34 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X267 VOUT.t228 pdrv1.t112 VDD.t258 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X268 VDD.t22 pdrv2.t84 VOUT.t21 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X269 vcomp VIN.t3 a_n551_n345# VDD.t452 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X270 VSS.t75 ndrv.t62 VOUT.t516 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X271 VOUT.t66 pdrv2.t85 VDD.t84 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X272 VDD.t463 pdrv2.t86 VOUT.t508 VDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X273 VDD.t257 pdrv1.t113 VOUT.t227 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X274 a_n3822_n3390# a_1610_n3072# VSS.t10 sky130_fd_pr__res_xhigh_po w=0.35 l=25
X275 VOUT.t226 pdrv1.t114 VDD.t256 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X276 VOUT.t501 pdrv2.t87 VDD.t456 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X277 VOUT.t14 ndrv.t63 VSS.t74 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X278 VOUT.t493 pdrv2.t88 VDD.t447 VDD.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X279 VDD.t123 pdrv2.t89 VOUT.t100 VDD.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X280 VDD.t255 pdrv1.t115 VOUT.t225 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X281 VDD.t250 pdrv1.t116 VOUT.t224 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X282 pdrv2 a_n3090_640# VDD.t60 VDD.t59 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X283 VDD.t254 pdrv1.t117 VOUT.t223 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X284 VDD.t253 pdrv1.t118 VOUT.t222 VDD.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X285 VDD.t252 pdrv1.t119 VOUT.t221 VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X286 VSS.t12 nbias.t2 nbias.t3 VSS.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X287 VOUT.t220 pdrv1.t120 VDD.t251 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X288 VOUT.t509 pdrv2.t90 VDD.t464 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X289 VOUT.t386 pdrv2.t91 VDD.t403 VDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X290 VDD.t389 pdrv2.t92 VOUT.t369 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
D0 VSS.t11 EN.t0 sky130_fd_pr__diode_pw2nd_05v5 pj=2.4e+06 area=3.6e+11
X291 VDD.t249 pdrv1.t121 VOUT.t219 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X292 VOUT.t218 pdrv1.t122 VDD.t248 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X293 VOUT.t346 ndrv.t64 VSS.t73 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X294 VOUT.t54 ndrv.t65 VSS.t72 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X295 VOUT.t217 pdrv1.t123 VDD.t247 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X296 VOUT.t133 pdrv2.t93 VDD.t166 VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X297 VOUT.t67 pdrv2.t94 VDD.t85 VDD.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X298 VOUT.t216 pdrv1.t124 VDD.t246 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X299 VDD.t148 pdrv2.t95 VOUT.t122 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X300 VDD.t245 pdrv1.t125 VOUT.t215 VDD.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X301 VOUT.t83 pdrv2.t96 VDD.t104 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X302 VOUT.t68 pdrv2.t97 VDD.t86 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X303 VOUT.t375 pdrv2.t98 VDD.t395 VDD.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X304 VDD.t49 pdrv2.t99 VOUT.t40 VDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X305 VOUT.t214 pdrv1.t126 VDD.t244 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X306 VDD.t167 pdrv2.t100 VOUT.t134 VDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X307 VOUT.t213 pdrv1.t127 VDD.t243 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X308 VDD.t396 pdrv2.t101 VOUT.t376 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X309 VOUT.t385 pdrv2.t102 VDD.t402 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X310 VSS.t71 ndrv.t66 VOUT.t511 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X311 VDD.t58 a_n3090_640# pdrv2 VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X312 VDD.t242 pdrv1.t128 VOUT.t212 VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X313 VOUT.t379 pdrv2.t103 VDD.t399 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X314 VDD.t5 pdrv2.t104 VOUT.t5 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X315 VDD.t241 pdrv1.t129 VOUT.t211 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X316 VDD.t457 pdrv2.t105 VOUT.t502 VDD.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X317 VOUT.t499 pdrv2.t106 VDD.t454 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X318 a_n1922_640# a_n1922_640# VDD.t156 VDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X319 VDD.t240 pdrv1.t130 VOUT.t210 VDD.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X320 VDD.t118 pdrv2.t107 VOUT.t95 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X321 VOUT.t387 ndrv.t67 VSS.t70 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X322 VOUT.t117 pdrv2.t108 VDD.t142 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X323 VSS.t69 ndrv.t68 VOUT.t55 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X324 VOUT.t378 pdrv2.t109 VDD.t398 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X325 VOUT.t344 pdrv2.t110 VDD.t372 VDD.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X326 VOUT.t209 pdrv1.t131 VDD.t239 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X327 VOUT.t490 pdrv2.t111 VDD.t443 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X328 vcomn2 nbias.t9 VSS.t8 VSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X329 VDD.t48 pdrv2.t112 VOUT.t39 VDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X330 VSS.t68 ndrv.t69 VOUT.t360 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X331 VOUT.t208 pdrv1.t132 VDD.t238 VDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X332 VDD.t237 pdrv1.t133 VOUT.t207 VDD.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X333 VDD.t147 pdrv2.t113 VOUT.t121 VDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X334 VOUT.t411 ndrv.t70 VSS.t67 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X335 VOUT.t471 ndrv.t71 VSS.t66 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X336 VDD.t236 pdrv1.t134 VOUT.t206 VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X337 VDD.t235 pdrv1.t135 VOUT.t205 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X338 VSS.t65 ndrv.t72 VOUT.t53 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X339 VOUT.t204 pdrv1.t136 VDD.t234 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X340 VOUT.t105 pdrv2.t114 VDD.t128 VDD.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X341 VOUT.t15 ndrv.t73 VSS.t64 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X342 VDD.t233 pdrv1.t137 VOUT.t203 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X343 VOUT.t367 pdrv2.t115 VDD.t387 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X344 VDD.t82 pdrv2.t116 VOUT.t65 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X345 VSS.t63 ndrv.t74 VOUT.t36 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X346 VSS.t62 ndrv.t75 VOUT.t362 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X347 VOUT.t202 pdrv1.t138 VDD.t232 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X348 VDD.t231 pdrv1.t139 VOUT.t201 VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X349 VDD.t230 pdrv1.t140 VOUT.t200 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X350 VOUT.t439 ndrv.t76 VSS.t61 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X351 VOUT.t199 pdrv1.t141 VDD.t229 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X352 vcomp VIP.t0 ndrv VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X353 VOUT.t124 pdrv2.t117 VDD.t150 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X354 VOUT.t96 pdrv2.t118 VDD.t119 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X355 VSS.t60 ndrv.t77 VOUT.t517 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X356 VOUT.t73 pdrv2.t119 VDD.t92 VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X357 VOUT.t64 pdrv2.t120 VDD.t81 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X358 VOUT.t198 pdrv1.t142 VDD.t228 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X359 VOUT.t512 pdrv2.t121 VDD.t465 VDD.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X360 VOUT.t500 pdrv2.t122 VDD.t455 VDD.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X361 a_n3822_n2754# a_1610_n3072# VSS.t14 sky130_fd_pr__res_xhigh_po w=0.35 l=25
X362 VDD.t227 pdrv1.t143 VOUT.t197 VDD.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X363 VDD.t94 pdrv2.t123 VOUT.t74 VDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X364 VOUT.t131 pdrv2.t124 VDD.t164 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X365 VDD.t226 pdrv1.t144 VOUT.t196 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X366 VSS.t59 ndrv.t78 VOUT.t396 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X367 VDD.t141 pdrv2.t125 VOUT.t116 VDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X368 pbias pbias VDD.t36 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X369 VOUT.t98 pdrv2.t126 VDD.t121 VDD.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X370 VOUT.t43 ndrv.t79 VSS.t58 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X371 VDD.t442 pdrv2.t127 VOUT.t489 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X372 VOUT.t432 ndrv.t80 VSS.t57 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X373 VDD.t225 pdrv1.t145 VOUT.t195 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X374 pdrv2 VIP.t1 vcomn2 VSS.t1 sky130_fd_pr__nfet_03v3_nvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X375 VOUT.t380 ndrv.t81 VSS.t56 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X376 VSS.t55 ndrv.t82 VOUT.t410 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X377 VDD.t391 pdrv2.t128 VOUT.t371 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X378 VOUT.t374 pdrv2.t129 VDD.t394 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X379 VSS.t54 ndrv.t83 VOUT.t442 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X380 VDD.t216 pdrv1.t146 VOUT.t194 VDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X381 VSS.t53 ndrv.t84 VOUT.t89 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X382 VDD.t224 pdrv1.t147 VOUT.t193 VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X383 VDD.t223 pdrv1.t148 VOUT.t192 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X384 VOUT.t341 ndrv.t85 VSS.t52 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X385 VDD.t163 pdrv2.t130 VOUT.t130 VDD.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X386 VOUT.t59 pdrv2.t131 VDD.t74 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X387 VDD.t222 pdrv1.t149 VOUT.t191 VDD.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X388 VOUT.t112 pdrv2.t132 VDD.t137 VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X389 VOUT.t465 ndrv.t86 VSS.t51 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X390 VDD.t56 a_n3090_640# a_n3090_640# VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X391 VOUT.t99 pdrv2.t133 VDD.t122 VDD.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X392 VDD.t32 pdrv2.t134 VOUT.t26 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X393 VOUT.t370 pdrv2.t135 VDD.t390 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X394 VOUT.t384 pdrv2.t136 VDD.t401 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X395 VOUT.t48 pdrv2.t137 VDD.t66 VDD.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X396 VDD.t215 pdrv1.t150 VOUT.t190 VDD.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X397 VOUT.t189 pdrv1.t151 VDD.t221 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X398 VSS.t50 ndrv.t87 VOUT.t392 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X399 VOUT.t188 pdrv1.t152 VDD.t220 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X400 VDD.t65 pdrv2.t138 VOUT.t47 VDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X401 VSS.t49 ndrv.t88 VOUT.t470 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X402 VOUT.t187 pdrv1.t153 VDD.t219 VDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X403 VSS.t48 ndrv.t89 VOUT.t347 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X404 VOUT.t186 pdrv1.t154 VDD.t218 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X405 VDD.t462 pdrv2.t139 VOUT.t507 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X406 VOUT.t400 ndrv.t90 VSS.t47 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X407 VDD.t103 pdrv2.t140 VOUT.t82 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X408 VOUT.t357 pdrv2.t141 VDD.t380 VDD.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X409 VOUT.t6 ndrv.t91 VSS.t46 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X410 VDD.t217 pdrv1.t155 VOUT.t185 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X411 VOUT.t184 pdrv1.t156 VDD.t214 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X412 VOUT.t348 ndrv.t92 VSS.t45 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X413 VDD.t453 pdrv2.t142 VOUT.t498 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X414 VSS.t138 nbias.t10 pbias VSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X415 VDD.t90 pdrv2.t143 VOUT.t72 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X416 VDD.t213 pdrv1.t157 VOUT.t183 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X417 VOUT.t94 pdrv2.t144 VDD.t116 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X418 VDD.t64 pdrv2.t145 VOUT.t46 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X419 VDD.t139 pdrv2.t146 VOUT.t115 VDD.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X420 VSS.t44 ndrv.t93 VOUT.t128 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X421 VSS.t43 ndrv.t94 VOUT.t481 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X422 VOUT.t4 pdrv2.t147 VDD.t3 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X423 VOUT.t182 pdrv1.t158 VDD.t212 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X424 VSS.t3 a_n551_n345# ndrv VSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X425 VOUT.t424 ndrv.t95 VSS.t42 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X426 VDD.t211 pdrv1.t159 VOUT.t181 VDD.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X427 VOUT.t486 pdrv2.t148 VDD.t439 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X428 VOUT.t497 pdrv2.t149 VDD.t451 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X429 VOUT.t519 ndrv.t96 VSS.t41 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X430 VOUT.t71 pdrv2.t150 VDD.t89 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X431 VDD.t62 pdrv2.t151 VOUT.t44 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X432 VOUT.t491 pdrv2.t152 VDD.t444 VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X433 VOUT.t63 pdrv2.t153 VDD.t79 VDD.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X434 VOUT.t119 pdrv2.t154 VDD.t145 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X435 VOUT.t31 ndrv.t97 VSS.t40 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X436 VOUT.t49 ndrv.t98 VSS.t39 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X437 VSS.t38 ndrv.t99 VOUT.t69 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X438 VSS.t37 ndrv.t100 VOUT.t113 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X439 pdrv1.t0 VIP.t2 vcomn1 VSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X440 VDD.t210 pdrv1.t160 VOUT.t180 VDD.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X441 VDD.t96 pdrv2.t155 VOUT.t76 VDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X442 VOUT.t179 pdrv1.t161 VDD.t209 VDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X443 VOUT.t354 ndrv.t101 VSS.t36 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X444 VDD.t208 pdrv1.t162 VOUT.t178 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X445 VSS.t35 ndrv.t102 VOUT.t510 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X446 VSS.t34 ndrv.t103 VOUT.t474 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X447 VDD.t100 pdrv2.t156 VOUT.t79 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X448 VOUT.t372 pdrv2.t157 VDD.t392 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X449 VOUT.t177 pdrv1.t163 VDD.t207 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X450 VOUT.t416 ndrv.t104 VSS.t33 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X451 VDD.t206 pdrv1.t164 VOUT.t176 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X452 VDD.t205 pdrv1.t165 VOUT.t175 VDD.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X453 VOUT.t174 pdrv1.t166 VDD.t204 VDD.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X454 VOUT.t488 pdrv2.t158 VDD.t441 VDD.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X455 VDD.t203 pdrv1.t167 VOUT.t173 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X456 VOUT.t28 ndrv.t105 VSS.t32 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X457 VSS.t31 ndrv.t106 VOUT.t345 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X458 VOUT.t420 ndrv.t107 VSS.t30 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X459 VDD.t202 pdrv1.t168 VOUT.t172 VDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X460 VSS.t29 ndrv.t108 VOUT.t30 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X461 VSS.t7 nbias.t0 nbias.t1 VSS.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X462 VDD.t201 pdrv1.t169 VOUT.t171 VDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X463 VDD.t99 pdrv2.t159 VOUT.t78 VDD.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X464 VOUT.t111 pdrv2.t160 VDD.t136 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X465 VOUT.t355 pdrv2.t161 VDD.t378 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X466 VOUT.t170 pdrv1.t170 VDD.t200 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X467 VSS.t28 ndrv.t109 VOUT.t479 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X468 VOUT.t169 pdrv1.t171 VDD.t199 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X469 VOUT.t473 ndrv.t110 VSS.t27 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X470 ndrv VIP.t3 vcomp VDD.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X471 VDD.t198 pdrv1.t172 VOUT.t168 VDD.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X472 VOUT.t92 pdrv2.t162 VDD.t113 VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X473 VOUT.t408 ndrv.t111 VSS.t26 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X474 VDD.t197 pdrv1.t173 VOUT.t167 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X475 VOUT.t81 pdrv2.t163 VDD.t102 VDD.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X476 VDD.t25 pdrv2.t164 VOUT.t22 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X477 VOUT.t166 pdrv1.t174 VDD.t191 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X478 VDD.t449 pdrv2.t165 VOUT.t495 VDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X479 VOUT.t61 pdrv2.t166 VDD.t75 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X480 VSS.t25 ndrv.t112 VOUT.t426 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X481 VSS.t24 ndrv.t113 VOUT.t7 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X482 VSS.t22 ndrv.t114 VOUT.t409 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X483 VDD.t196 pdrv1.t175 VOUT.t165 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X484 VDD.t195 pdrv1.t176 VOUT.t164 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X485 VDD.t149 pdrv2.t167 VOUT.t123 VDD.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X486 VOUT.t163 pdrv1.t177 VDD.t194 VDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X487 VOUT.t162 pdrv1.t178 VDD.t193 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X488 VDD.t30 pdrv2.t168 VOUT.t25 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X489 a_1610_n2436# EN.t1 nbias.t8 VSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X490 VSS.t21 ndrv.t115 VOUT.t359 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X491 VDD.t146 pdrv2.t169 VOUT.t120 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X492 VDD.t134 pdrv2.t170 VOUT.t110 VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X493 VDD.t192 pdrv1.t179 VOUT.t161 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X494 vcomn1 nbias.t11 VSS.t13 VSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X495 VOUT.t160 pdrv1.t180 VDD.t190 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X496 VSS.t20 ndrv.t116 VOUT.t417 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X497 VDD.t138 pdrv2.t171 VOUT.t114 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X498 a_n3822_n2754# a_1610_n2436# VSS.t0 sky130_fd_pr__res_xhigh_po w=0.35 l=25
X499 VDD.t28 pdrv2.t172 VOUT.t24 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X500 VDD.t189 pdrv1.t181 VOUT.t159 VDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X501 VOUT.t356 pdrv2.t173 VDD.t379 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X502 VDD.t382 pdrv2.t174 VOUT.t361 VDD.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X503 VOUT.t390 pdrv2.t175 VDD.t406 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X504 VOUT.t158 pdrv1.t182 VDD.t186 VDD.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X505 VDD.t188 pdrv1.t183 VOUT.t157 VDD.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X506 VOUT.t506 pdrv2.t176 VDD.t461 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X507 VDD.t385 pdrv2.t177 VOUT.t365 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X508 a_n3090_640# a_n3090_640# VDD.t54 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X509 VOUT.t156 pdrv1.t184 VDD.t185 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X510 VOUT.t77 pdrv2.t178 VDD.t97 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X511 VOUT.t407 ndrv.t117 VSS.t19 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X512 VOUT.t388 pdrv2.t179 VDD.t404 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X513 VDD.t440 pdrv2.t180 VOUT.t487 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X514 VOUT.t366 pdrv2.t181 VDD.t386 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X515 VOUT.t23 pdrv2.t182 VDD.t26 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X516 VDD.t405 pdrv2.t183 VOUT.t389 VDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X517 VSS.t18 ndrv.t118 VOUT.t33 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X518 VDD.t101 pdrv2.t184 VOUT.t80 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X519 VOUT.t431 ndrv.t119 VSS.t16 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X520 VOUT.t155 pdrv1.t185 VDD.t181 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X521 VOUT.t154 pdrv1.t186 VDD.t184 VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X522 VDD.t183 pdrv1.t187 VOUT.t153 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X523 VOUT.t152 pdrv1.t188 VDD.t182 VDD.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X524 VOUT.t62 pdrv2.t185 VDD.t77 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X525 VOUT.t151 pdrv1.t189 VDD.t180 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X526 VDD.t20 pdrv2.t186 VOUT.t20 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X527 VOUT.t150 pdrv1.t190 VDD.t179 VDD.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X528 VDD.t384 pdrv2.t187 VOUT.t364 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X529 VOUT.t149 pdrv1.t191 VDD.t178 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X530 VDD.t177 pdrv1.t192 VOUT.t148 VDD.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X531 VDD.t176 pdrv1.t193 VOUT.t147 VDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X532 VDD.t175 pdrv1.t194 VOUT.t146 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X533 VDD.t174 pdrv1.t195 VOUT.t145 VDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X534 VOUT.t58 pdrv2.t188 VDD.t73 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X535 VOUT.t492 pdrv2.t189 VDD.t445 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X536 VDD.t450 pdrv2.t190 VOUT.t496 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X537 VOUT.t505 pdrv2.t191 VDD.t460 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X538 VDD.t63 pdrv2.t192 VOUT.t45 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X539 VOUT.t373 pdrv2.t193 VDD.t393 VDD.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X540 VOUT.t144 pdrv1.t196 VDD.t173 VDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X541 VOUT.t57 pdrv2.t194 VDD.t71 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X542 VDD.t172 pdrv1.t197 VOUT.t143 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X543 VOUT.t142 pdrv1.t198 VDD.t171 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X544 VDD.t114 pdrv2.t195 VOUT.t93 VDD.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X545 VDD.t170 pdrv1.t199 VOUT.t141 VDD.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X546 VOUT.t140 pdrv1.t200 VDD.t169 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X547 VOUT.t3 pdrv2.t196 VDD.t1 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X548 a_n3822_n3390# VDD.t23 VSS.t2 sky130_fd_pr__res_xhigh_po w=0.35 l=25
X549 VDD.t168 pdrv1.t201 VOUT.t139 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X550 VOUT.t504 pdrv2.t197 VDD.t459 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X551 VDD.t144 pdrv2.t198 VOUT.t118 VDD.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
X552 VDD.t458 pdrv2.t199 VOUT.t503 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.5
R0 pdrv1.n37 pdrv1.t118 92.48
R1 pdrv1.n38 pdrv1.t17 92.48
R2 pdrv1.n38 pdrv1.t23 92.48
R3 pdrv1.n39 pdrv1.t136 92.48
R4 pdrv1.n39 pdrv1.t96 92.48
R5 pdrv1.n40 pdrv1.t47 92.48
R6 pdrv1.n40 pdrv1.t147 92.48
R7 pdrv1.n41 pdrv1.t100 92.48
R8 pdrv1.n41 pdrv1.t19 92.48
R9 pdrv1.n42 pdrv1.t69 92.48
R10 pdrv1.n42 pdrv1.t119 92.48
R11 pdrv1.n43 pdrv1.t2 92.48
R12 pdrv1.n43 pdrv1.t195 92.48
R13 pdrv1.n44 pdrv1.t103 92.48
R14 pdrv1.n44 pdrv1.t148 92.48
R15 pdrv1.n45 pdrv1.t48 92.48
R16 pdrv1.n45 pdrv1.t97 92.48
R17 pdrv1.n46 pdrv1.t89 92.48
R18 pdrv1.n46 pdrv1.t172 92.48
R19 pdrv1.n47 pdrv1.t18 92.48
R20 pdrv1.n47 pdrv1.t179 92.48
R21 pdrv1.n48 pdrv1.t24 92.48
R22 pdrv1.n48 pdrv1.t77 92.48
R23 pdrv1.n49 pdrv1.t124 92.48
R24 pdrv1.n49 pdrv1.t157 92.48
R25 pdrv1.n50 pdrv1.t56 92.48
R26 pdrv1.n50 pdrv1.t160 92.48
R27 pdrv1.n51 pdrv1.t6 92.48
R28 pdrv1.n51 pdrv1.t54 92.48
R29 pdrv1.n52 pdrv1.t105 92.48
R30 pdrv1.n52 pdrv1.t187 92.48
R31 pdrv1.n53 pdrv1.t34 92.48
R32 pdrv1.n53 pdrv1.t87 92.48
R33 pdrv1.n19 pdrv1.t5 92.4691
R34 pdrv1.n19 pdrv1.t121 92.4691
R35 pdrv1.n19 pdrv1.t196 92.4691
R36 pdrv1.n19 pdrv1.t113 92.4691
R37 pdrv1.n18 pdrv1.t122 92.4691
R38 pdrv1.n18 pdrv1.t76 92.4691
R39 pdrv1.n18 pdrv1.t171 92.4691
R40 pdrv1.n18 pdrv1.t133 92.4691
R41 pdrv1.n17 pdrv1.t39 92.4691
R42 pdrv1.n17 pdrv1.t51 92.4691
R43 pdrv1.n17 pdrv1.t151 92.4691
R44 pdrv1.n17 pdrv1.t116 92.4691
R45 pdrv1.n16 pdrv1.t67 92.4691
R46 pdrv1.n16 pdrv1.t165 92.4691
R47 pdrv1.n16 pdrv1.t120 92.4691
R48 pdrv1.n16 pdrv1.t46 92.4691
R49 pdrv1.n15 pdrv1.t95 92.4691
R50 pdrv1.n15 pdrv1.t134 92.4691
R51 pdrv1.n15 pdrv1.t22 92.4691
R52 pdrv1.n15 pdrv1.t15 92.4691
R53 pdrv1.n14 pdrv1.t123 92.4691
R54 pdrv1.n14 pdrv1.t167 92.4691
R55 pdrv1.n14 pdrv1.t68 92.4691
R56 pdrv1.n14 pdrv1.t117 92.4691
R57 pdrv1.n13 pdrv1.t111 92.4691
R58 pdrv1.n13 pdrv1.t192 92.4691
R59 pdrv1.n13 pdrv1.t40 92.4691
R60 pdrv1.n13 pdrv1.t201 92.4691
R61 pdrv1.n12 pdrv1.t52 92.4691
R62 pdrv1.n12 pdrv1.t99 92.4691
R63 pdrv1.n12 pdrv1.t138 92.4691
R64 pdrv1.n12 pdrv1.t176 92.4691
R65 pdrv1.n11 pdrv1.t82 92.4691
R66 pdrv1.n11 pdrv1.t183 92.4691
R67 pdrv1.n11 pdrv1.t28 92.4691
R68 pdrv1.n11 pdrv1.t80 92.4691
R69 pdrv1.n10 pdrv1.t126 92.4691
R70 pdrv1.n10 pdrv1.t9 92.4691
R71 pdrv1.n10 pdrv1.t60 92.4691
R72 pdrv1.n10 pdrv1.t109 92.4691
R73 pdrv1.n20 pdrv1.t27 92.4664
R74 pdrv1.n20 pdrv1.t182 92.4664
R75 pdrv1.n20 pdrv1.t144 92.4664
R76 pdrv1.n20 pdrv1.t50 92.4664
R77 pdrv1.n21 pdrv1.t199 92.4664
R78 pdrv1.n21 pdrv1.t156 92.4664
R79 pdrv1.n21 pdrv1.t125 92.4664
R80 pdrv1.n21 pdrv1.t200 92.4664
R81 pdrv1.n22 pdrv1.t115 92.4664
R82 pdrv1.n22 pdrv1.t66 92.4664
R83 pdrv1.n22 pdrv1.t16 92.4664
R84 pdrv1.n22 pdrv1.t174 92.4664
R85 pdrv1.n23 pdrv1.t135 92.4664
R86 pdrv1.n23 pdrv1.t166 92.4664
R87 pdrv1.n23 pdrv1.t130 92.4664
R88 pdrv1.n23 pdrv1.t30 92.4664
R89 pdrv1.n24 pdrv1.t36 92.4664
R90 pdrv1.n24 pdrv1.t188 92.4664
R91 pdrv1.n24 pdrv1.t108 92.4664
R92 pdrv1.n24 pdrv1.t45 92.4664
R93 pdrv1.n25 pdrv1.t146 92.4664
R94 pdrv1.n25 pdrv1.t154 92.4664
R95 pdrv1.n25 pdrv1.t63 92.4664
R96 pdrv1.n25 pdrv1.t12 92.4664
R97 pdrv1.n26 pdrv1.t168 92.4664
R98 pdrv1.n26 pdrv1.t41 92.4664
R99 pdrv1.n26 pdrv1.t107 92.4664
R100 pdrv1.n26 pdrv1.t186 92.4664
R101 pdrv1.n27 pdrv1.t35 92.4664
R102 pdrv1.n27 pdrv1.t90 92.4664
R103 pdrv1.n27 pdrv1.t173 92.4664
R104 pdrv1.n27 pdrv1.t163 92.4664
R105 pdrv1.n28 pdrv1.t61 92.4664
R106 pdrv1.n28 pdrv1.t112 92.4664
R107 pdrv1.n28 pdrv1.t194 92.4664
R108 pdrv1.n28 pdrv1.t44 92.4664
R109 pdrv1.n29 pdrv1.t33 92.4664
R110 pdrv1.n29 pdrv1.t132 92.4664
R111 pdrv1.n29 pdrv1.t43 92.4664
R112 pdrv1.n29 pdrv1.t141 92.4664
R113 pdrv1.n9 pdrv1.t158 92.4637
R114 pdrv1.n9 pdrv1.t72 92.4637
R115 pdrv1.n9 pdrv1.t153 92.4637
R116 pdrv1.n9 pdrv1.t62 92.4637
R117 pdrv1.n8 pdrv1.t74 92.4637
R118 pdrv1.n8 pdrv1.t20 92.4637
R119 pdrv1.n8 pdrv1.t131 92.4637
R120 pdrv1.n8 pdrv1.t91 92.4637
R121 pdrv1.n7 pdrv1.t189 92.4637
R122 pdrv1.n7 pdrv1.t197 92.4637
R123 pdrv1.n7 pdrv1.t114 92.4637
R124 pdrv1.n7 pdrv1.t64 92.4637
R125 pdrv1.n6 pdrv1.t13 92.4637
R126 pdrv1.n6 pdrv1.t128 92.4637
R127 pdrv1.n6 pdrv1.t71 92.4637
R128 pdrv1.n6 pdrv1.t193 92.4637
R129 pdrv1.n5 pdrv1.t42 92.4637
R130 pdrv1.n5 pdrv1.t94 92.4637
R131 pdrv1.n5 pdrv1.t178 92.4637
R132 pdrv1.n5 pdrv1.t169 92.4637
R133 pdrv1.n4 pdrv1.t75 92.4637
R134 pdrv1.n4 pdrv1.t129 92.4637
R135 pdrv1.n4 pdrv1.t14 92.4637
R136 pdrv1.n4 pdrv1.t65 92.4637
R137 pdrv1.n3 pdrv1.t58 92.4637
R138 pdrv1.n3 pdrv1.t149 92.4637
R139 pdrv1.n3 pdrv1.t190 92.4637
R140 pdrv1.n3 pdrv1.t155 92.4637
R141 pdrv1.n2 pdrv1.t198 92.4637
R142 pdrv1.n2 pdrv1.t49 92.4637
R143 pdrv1.n2 pdrv1.t98 92.4637
R144 pdrv1.n2 pdrv1.t137 92.4637
R145 pdrv1.n1 pdrv1.t26 92.4637
R146 pdrv1.n1 pdrv1.t143 92.4637
R147 pdrv1.n1 pdrv1.t180 92.4637
R148 pdrv1.n1 pdrv1.t25 92.4637
R149 pdrv1.n0 pdrv1.t79 92.4637
R150 pdrv1.n0 pdrv1.t162 92.4637
R151 pdrv1.n0 pdrv1.t8 92.4637
R152 pdrv1.n0 pdrv1.t57 92.4637
R153 pdrv1.n33 pdrv1.t184 92.4623
R154 pdrv1.n35 pdrv1.t170 92.4623
R155 pdrv1.n33 pdrv1.t101 92.4623
R156 pdrv1.n35 pdrv1.t85 92.4623
R157 pdrv1.n32 pdrv1.t177 92.4623
R158 pdrv1.n34 pdrv1.t161 92.4623
R159 pdrv1.n32 pdrv1.t93 92.4623
R160 pdrv1.n34 pdrv1.t78 92.4623
R161 pdrv1.n31 pdrv1.t102 92.4623
R162 pdrv1.n36 pdrv1.t86 92.4623
R163 pdrv1.n31 pdrv1.t53 92.4623
R164 pdrv1.n36 pdrv1.t32 92.4623
R165 pdrv1.n30 pdrv1.t152 92.4623
R166 pdrv1.n37 pdrv1.t142 92.4623
R167 pdrv1.n37 pdrv1.t104 92.4623
R168 pdrv1.n38 pdrv1.t3 92.4623
R169 pdrv1.n38 pdrv1.t10 92.4623
R170 pdrv1.n39 pdrv1.t127 92.4623
R171 pdrv1.n39 pdrv1.t81 92.4623
R172 pdrv1.n40 pdrv1.t29 92.4623
R173 pdrv1.n40 pdrv1.t139 92.4623
R174 pdrv1.n41 pdrv1.t84 92.4623
R175 pdrv1.n41 pdrv1.t7 92.4623
R176 pdrv1.n42 pdrv1.t55 92.4623
R177 pdrv1.n5 pdrv1.t106 92.4623
R178 pdrv1.n5 pdrv1.t185 92.4623
R179 pdrv1.n5 pdrv1.t181 92.4623
R180 pdrv1.n4 pdrv1.t88 92.4623
R181 pdrv1.n4 pdrv1.t140 92.4623
R182 pdrv1.n4 pdrv1.t31 92.4623
R183 pdrv1.n4 pdrv1.t83 92.4623
R184 pdrv1.n3 pdrv1.t73 92.4623
R185 pdrv1.n3 pdrv1.t159 92.4623
R186 pdrv1.n3 pdrv1.t4 92.4623
R187 pdrv1.n3 pdrv1.t164 92.4623
R188 pdrv1.n2 pdrv1.t11 92.4623
R189 pdrv1.n2 pdrv1.t59 92.4623
R190 pdrv1.n2 pdrv1.t110 92.4623
R191 pdrv1.n2 pdrv1.t145 92.4623
R192 pdrv1.n1 pdrv1.t38 92.4623
R193 pdrv1.n1 pdrv1.t150 92.4623
R194 pdrv1.n1 pdrv1.t191 92.4623
R195 pdrv1.n1 pdrv1.t37 92.4623
R196 pdrv1.n0 pdrv1.t92 92.4623
R197 pdrv1.n0 pdrv1.t175 92.4623
R198 pdrv1.n0 pdrv1.t21 92.4623
R199 pdrv1.n0 pdrv1.t70 92.4623
R200 pdrv1.t1 pdrv1.t0 23.7687
R201 pdrv1.n30 pdrv1.n57 8.59371
R202 pdrv1 pdrv1.t1 7.33433
R203 pdrv1 pdrv1.n58 4.80282
R204 pdrv1.n58 pdrv1.n56 0.639172
R205 pdrv1.n56 pdrv1.n55 0.6255
R206 pdrv1.n55 pdrv1.n54 0.619641
R207 pdrv1.n33 pdrv1.n32 0.573381
R208 pdrv1.n32 pdrv1.n31 0.573381
R209 pdrv1.n31 pdrv1.n30 0.573381
R210 pdrv1.n56 pdrv1.n35 0.487342
R211 pdrv1.n52 pdrv1.n53 0.416289
R212 pdrv1.n51 pdrv1.n52 0.416289
R213 pdrv1.n50 pdrv1.n51 0.416289
R214 pdrv1.n49 pdrv1.n50 0.416289
R215 pdrv1.n48 pdrv1.n49 0.416289
R216 pdrv1.n47 pdrv1.n48 0.416289
R217 pdrv1.n46 pdrv1.n47 0.416289
R218 pdrv1.n45 pdrv1.n46 0.416289
R219 pdrv1.n44 pdrv1.n45 0.416289
R220 pdrv1.n43 pdrv1.n44 0.416289
R221 pdrv1.n42 pdrv1.n43 0.416289
R222 pdrv1.n41 pdrv1.n42 0.416289
R223 pdrv1.n40 pdrv1.n41 0.416289
R224 pdrv1.n39 pdrv1.n40 0.416289
R225 pdrv1.n38 pdrv1.n39 0.416289
R226 pdrv1.n37 pdrv1.n38 0.416289
R227 pdrv1.n36 pdrv1.n37 0.416289
R228 pdrv1.n34 pdrv1.n36 0.416289
R229 pdrv1.n35 pdrv1.n34 0.416289
R230 pdrv1.n58 pdrv1.n33 0.403486
R231 pdrv1.n55 pdrv1.n9 0.402674
R232 pdrv1.n54 pdrv1.n19 0.402674
R233 pdrv1.n54 pdrv1.n29 1.03353
R234 pdrv1.n21 pdrv1.n20 1.03093
R235 pdrv1.n11 pdrv1.n10 1.03093
R236 pdrv1.n1 pdrv1.n0 1.03093
R237 pdrv1.n29 pdrv1.n28 0.687457
R238 pdrv1.n28 pdrv1.n27 0.687457
R239 pdrv1.n27 pdrv1.n26 0.687457
R240 pdrv1.n26 pdrv1.n25 0.687457
R241 pdrv1.n25 pdrv1.n24 0.687457
R242 pdrv1.n24 pdrv1.n23 0.687457
R243 pdrv1.n23 pdrv1.n22 0.687457
R244 pdrv1.n22 pdrv1.n21 0.687457
R245 pdrv1.n19 pdrv1.n18 0.687457
R246 pdrv1.n18 pdrv1.n17 0.687457
R247 pdrv1.n17 pdrv1.n16 0.687457
R248 pdrv1.n16 pdrv1.n15 0.687457
R249 pdrv1.n15 pdrv1.n14 0.687457
R250 pdrv1.n14 pdrv1.n13 0.687457
R251 pdrv1.n13 pdrv1.n12 0.687457
R252 pdrv1.n12 pdrv1.n11 0.687457
R253 pdrv1.n9 pdrv1.n8 0.687457
R254 pdrv1.n8 pdrv1.n7 0.687457
R255 pdrv1.n7 pdrv1.n6 0.687457
R256 pdrv1.n6 pdrv1.n5 0.687457
R257 pdrv1.n5 pdrv1.n4 0.687457
R258 pdrv1.n4 pdrv1.n3 0.687457
R259 pdrv1.n3 pdrv1.n2 0.687457
R260 pdrv1.n2 pdrv1.n1 0.687457
R261 VDD.n2996 VDD.n2835 190.655
R262 VDD.n5264 VDD.n5155 178.863
R263 VDD.n1251 VDD.n1247 133.655
R264 VDD.n1236 VDD.n1235 133.655
R265 VDD.n1708 VDD.n1704 133.655
R266 VDD.n1693 VDD.n1692 133.655
R267 VDD.n1686 VDD.n1682 133.655
R268 VDD.n1671 VDD.n1670 133.655
R269 VDD.n1552 VDD.n1548 133.655
R270 VDD.n1537 VDD.n1536 133.655
R271 VDD.n1570 VDD.n1566 133.655
R272 VDD.n1555 VDD.n1554 133.655
R273 VDD.n1233 VDD.n1229 133.655
R274 VDD.n1324 VDD.n1323 133.655
R275 VDD.n1444 VDD.n1440 133.655
R276 VDD.n1380 VDD.n1379 133.655
R277 VDD.n2781 VDD.n2780 92.5005
R278 VDD.n2778 VDD.n2777 92.5005
R279 VDD.n2775 VDD.n2774 92.5005
R280 VDD.n2772 VDD.n2771 92.5005
R281 VDD.n2769 VDD.n2768 92.5005
R282 VDD.n2766 VDD.n2765 92.5005
R283 VDD.n2763 VDD.n2762 92.5005
R284 VDD.n2760 VDD.n2759 92.5005
R285 VDD.n2757 VDD.n2756 92.5005
R286 VDD.n2754 VDD.n2753 92.5005
R287 VDD.n2751 VDD.n2750 92.5005
R288 VDD.n2748 VDD.n2747 92.5005
R289 VDD.n2745 VDD.n2744 92.5005
R290 VDD.n2742 VDD.n2741 92.5005
R291 VDD.n2739 VDD.n2738 92.5005
R292 VDD.n2736 VDD.n2735 92.5005
R293 VDD.n2733 VDD.n2732 92.5005
R294 VDD.n2787 VDD.n2786 92.5005
R295 VDD.n2785 VDD.n2784 92.5005
R296 VDD.n1080 VDD.n1079 92.5005
R297 VDD.n1076 VDD.n1075 92.5005
R298 VDD.n1072 VDD.n1071 92.5005
R299 VDD.n1068 VDD.n1067 92.5005
R300 VDD.n1064 VDD.n1063 92.5005
R301 VDD.n1060 VDD.n1059 92.5005
R302 VDD.n1056 VDD.n1055 92.5005
R303 VDD.n1053 VDD.n1052 92.5005
R304 VDD.n1050 VDD.n1049 92.5005
R305 VDD.n1047 VDD.n1046 92.5005
R306 VDD.n1044 VDD.n1043 92.5005
R307 VDD.n1041 VDD.n1040 92.5005
R308 VDD.n1038 VDD.n1037 92.5005
R309 VDD.n1035 VDD.n1034 92.5005
R310 VDD.n1032 VDD.n1031 92.5005
R311 VDD.n1029 VDD.n1028 92.5005
R312 VDD.n1026 VDD.n1025 92.5005
R313 VDD.n1023 VDD.n1022 92.5005
R314 VDD.n1020 VDD.n1019 92.5005
R315 VDD.n2790 VDD.n2789 92.5005
R316 VDD.n2793 VDD.n2792 92.5005
R317 VDD.n2796 VDD.n2795 92.5005
R318 VDD.n2799 VDD.n2798 92.5005
R319 VDD.n2802 VDD.n2801 92.5005
R320 VDD.n2805 VDD.n2804 92.5005
R321 VDD.n2808 VDD.n2807 92.5005
R322 VDD.n2811 VDD.n2810 92.5005
R323 VDD.n2814 VDD.n2813 92.5005
R324 VDD.n2817 VDD.n2816 92.5005
R325 VDD.n2820 VDD.n2819 92.5005
R326 VDD.n2823 VDD.n2822 92.5005
R327 VDD.n2826 VDD.n2825 92.5005
R328 VDD.n2830 VDD.n2829 92.5005
R329 VDD.n2832 VDD.n2831 92.5005
R330 VDD.n2894 VDD.n2893 92.5005
R331 VDD.n2896 VDD.n2895 92.5005
R332 VDD.n2898 VDD.n2897 92.5005
R333 VDD.n2989 VDD.n2988 92.5005
R334 VDD.n2991 VDD.n2990 92.5005
R335 VDD.n3031 VDD.n3030 92.5005
R336 VDD.n3010 VDD.n3009 92.5005
R337 VDD.n3395 VDD.n3394 92.5005
R338 VDD.n3415 VDD.n3414 92.5005
R339 VDD.n3436 VDD.n3435 92.5005
R340 VDD.n3456 VDD.n3455 92.5005
R341 VDD.n3477 VDD.n3476 92.5005
R342 VDD.n3500 VDD.n3499 92.5005
R343 VDD.n3507 VDD.n3506 92.5005
R344 VDD.n3544 VDD.n3543 92.5005
R345 VDD.n3548 VDD.n3547 92.5005
R346 VDD.n3567 VDD.n3566 92.5005
R347 VDD.n3587 VDD.n3586 92.5005
R348 VDD.n3608 VDD.n3607 92.5005
R349 VDD.n3626 VDD.n3625 92.5005
R350 VDD.n3650 VDD.n3649 92.5005
R351 VDD.n3674 VDD.n3673 92.5005
R352 VDD.n3697 VDD.n3696 92.5005
R353 VDD.n3718 VDD.n3717 92.5005
R354 VDD.n3737 VDD.n3736 92.5005
R355 VDD.n3757 VDD.n3756 92.5005
R356 VDD.n3777 VDD.n3776 92.5005
R357 VDD.n3797 VDD.n3796 92.5005
R358 VDD.n3818 VDD.n3817 92.5005
R359 VDD.n3841 VDD.n3840 92.5005
R360 VDD.n3864 VDD.n3863 92.5005
R361 VDD.n3873 VDD.n3872 92.5005
R362 VDD.n3869 VDD.n3868 92.5005
R363 VDD.n3909 VDD.n3908 92.5005
R364 VDD.n3926 VDD.n3925 92.5005
R365 VDD.n3947 VDD.n3946 92.5005
R366 VDD.n3965 VDD.n3964 92.5005
R367 VDD.n3990 VDD.n3989 92.5005
R368 VDD.n4014 VDD.n4013 92.5005
R369 VDD.n6574 VDD.n6573 92.5005
R370 VDD.n6577 VDD.n6576 92.5005
R371 VDD.n6581 VDD.n6580 92.5005
R372 VDD.n6585 VDD.n6584 92.5005
R373 VDD.n6589 VDD.n6588 92.5005
R374 VDD.n6593 VDD.n6592 92.5005
R375 VDD.n6597 VDD.n6596 92.5005
R376 VDD.n6601 VDD.n6600 92.5005
R377 VDD.n6605 VDD.n6604 92.5005
R378 VDD.n6609 VDD.n6608 92.5005
R379 VDD.n6613 VDD.n6612 92.5005
R380 VDD.n6617 VDD.n6616 92.5005
R381 VDD.n6621 VDD.n6620 92.5005
R382 VDD.n6693 VDD.n6692 92.5005
R383 VDD.n6689 VDD.n6688 92.5005
R384 VDD.n6685 VDD.n6684 92.5005
R385 VDD.n6681 VDD.n6680 92.5005
R386 VDD.n6677 VDD.n6676 92.5005
R387 VDD.n6673 VDD.n6672 92.5005
R388 VDD.n6669 VDD.n6668 92.5005
R389 VDD.n6665 VDD.n6664 92.5005
R390 VDD.n6661 VDD.n6660 92.5005
R391 VDD.n6657 VDD.n6656 92.5005
R392 VDD.n6653 VDD.n6652 92.5005
R393 VDD.n4470 VDD.n4469 92.5005
R394 VDD.n4494 VDD.n4493 92.5005
R395 VDD.n4516 VDD.n4515 92.5005
R396 VDD.n4521 VDD.n4520 92.5005
R397 VDD.n4541 VDD.n4540 92.5005
R398 VDD.n4571 VDD.n4570 92.5005
R399 VDD.n4575 VDD.n4574 92.5005
R400 VDD.n4593 VDD.n4592 92.5005
R401 VDD.n4617 VDD.n4616 92.5005
R402 VDD.n4640 VDD.n4639 92.5005
R403 VDD.n4663 VDD.n4662 92.5005
R404 VDD.n4685 VDD.n4684 92.5005
R405 VDD.n4704 VDD.n4703 92.5005
R406 VDD.n4724 VDD.n4723 92.5005
R407 VDD.n4743 VDD.n4742 92.5005
R408 VDD.n4762 VDD.n4761 92.5005
R409 VDD.n4779 VDD.n4778 92.5005
R410 VDD.n4802 VDD.n4801 92.5005
R411 VDD.n4826 VDD.n4825 92.5005
R412 VDD.n4831 VDD.n4830 92.5005
R413 VDD.n4868 VDD.n4867 92.5005
R414 VDD.n4888 VDD.n4887 92.5005
R415 VDD.n4895 VDD.n4894 92.5005
R416 VDD.n4927 VDD.n4926 92.5005
R417 VDD.n4931 VDD.n4930 92.5005
R418 VDD.n4951 VDD.n4950 92.5005
R419 VDD.n4974 VDD.n4973 92.5005
R420 VDD.n4998 VDD.n4997 92.5005
R421 VDD.n5019 VDD.n5018 92.5005
R422 VDD.n5038 VDD.n5037 92.5005
R423 VDD.n5058 VDD.n5057 92.5005
R424 VDD.n6466 VDD.n6465 92.5005
R425 VDD.n6469 VDD.n6468 92.5005
R426 VDD.n6473 VDD.n6472 92.5005
R427 VDD.n6477 VDD.n6476 92.5005
R428 VDD.n6481 VDD.n6480 92.5005
R429 VDD.n6485 VDD.n6484 92.5005
R430 VDD.n2994 VDD.n2993 92.5005
R431 VDD.n3034 VDD.n3033 92.5005
R432 VDD.n3013 VDD.n3012 92.5005
R433 VDD.n3398 VDD.n3397 92.5005
R434 VDD.n3418 VDD.n3417 92.5005
R435 VDD.n3439 VDD.n3438 92.5005
R436 VDD.n3459 VDD.n3458 92.5005
R437 VDD.n3480 VDD.n3479 92.5005
R438 VDD.n3503 VDD.n3502 92.5005
R439 VDD.n3505 VDD.n3504 92.5005
R440 VDD.n3546 VDD.n3545 92.5005
R441 VDD.n3551 VDD.n3550 92.5005
R442 VDD.n3570 VDD.n3569 92.5005
R443 VDD.n3590 VDD.n3589 92.5005
R444 VDD.n3611 VDD.n3610 92.5005
R445 VDD.n3629 VDD.n3628 92.5005
R446 VDD.n3653 VDD.n3652 92.5005
R447 VDD.n3677 VDD.n3676 92.5005
R448 VDD.n3700 VDD.n3699 92.5005
R449 VDD.n3721 VDD.n3720 92.5005
R450 VDD.n3740 VDD.n3739 92.5005
R451 VDD.n3760 VDD.n3759 92.5005
R452 VDD.n3780 VDD.n3779 92.5005
R453 VDD.n3800 VDD.n3799 92.5005
R454 VDD.n3821 VDD.n3820 92.5005
R455 VDD.n3844 VDD.n3843 92.5005
R456 VDD.n3867 VDD.n3866 92.5005
R457 VDD.n3871 VDD.n3870 92.5005
R458 VDD.n3907 VDD.n3906 92.5005
R459 VDD.n3912 VDD.n3911 92.5005
R460 VDD.n3929 VDD.n3928 92.5005
R461 VDD.n3950 VDD.n3949 92.5005
R462 VDD.n3968 VDD.n3967 92.5005
R463 VDD.n3993 VDD.n3992 92.5005
R464 VDD.n4017 VDD.n4016 92.5005
R465 VDD.n4039 VDD.n4038 92.5005
R466 VDD.n6579 VDD.n6578 92.5005
R467 VDD.n6583 VDD.n6582 92.5005
R468 VDD.n6587 VDD.n6586 92.5005
R469 VDD.n6591 VDD.n6590 92.5005
R470 VDD.n6595 VDD.n6594 92.5005
R471 VDD.n6599 VDD.n6598 92.5005
R472 VDD.n6603 VDD.n6602 92.5005
R473 VDD.n6607 VDD.n6606 92.5005
R474 VDD.n6611 VDD.n6610 92.5005
R475 VDD.n6615 VDD.n6614 92.5005
R476 VDD.n6619 VDD.n6618 92.5005
R477 VDD.n6695 VDD.n6694 92.5005
R478 VDD.n6691 VDD.n6690 92.5005
R479 VDD.n6687 VDD.n6686 92.5005
R480 VDD.n6683 VDD.n6682 92.5005
R481 VDD.n6679 VDD.n6678 92.5005
R482 VDD.n6675 VDD.n6674 92.5005
R483 VDD.n6671 VDD.n6670 92.5005
R484 VDD.n6667 VDD.n6666 92.5005
R485 VDD.n6663 VDD.n6662 92.5005
R486 VDD.n6659 VDD.n6658 92.5005
R487 VDD.n6655 VDD.n6654 92.5005
R488 VDD.n4452 VDD.n4451 92.5005
R489 VDD.n4473 VDD.n4472 92.5005
R490 VDD.n4497 VDD.n4496 92.5005
R491 VDD.n4519 VDD.n4518 92.5005
R492 VDD.n4537 VDD.n4536 92.5005
R493 VDD.n4539 VDD.n4538 92.5005
R494 VDD.n4573 VDD.n4572 92.5005
R495 VDD.n4578 VDD.n4577 92.5005
R496 VDD.n4596 VDD.n4595 92.5005
R497 VDD.n4620 VDD.n4619 92.5005
R498 VDD.n4643 VDD.n4642 92.5005
R499 VDD.n4666 VDD.n4665 92.5005
R500 VDD.n4688 VDD.n4687 92.5005
R501 VDD.n4707 VDD.n4706 92.5005
R502 VDD.n4727 VDD.n4726 92.5005
R503 VDD.n4746 VDD.n4745 92.5005
R504 VDD.n4765 VDD.n4764 92.5005
R505 VDD.n4782 VDD.n4781 92.5005
R506 VDD.n4805 VDD.n4804 92.5005
R507 VDD.n4829 VDD.n4828 92.5005
R508 VDD.n4852 VDD.n4851 92.5005
R509 VDD.n4871 VDD.n4870 92.5005
R510 VDD.n4891 VDD.n4890 92.5005
R511 VDD.n4893 VDD.n4892 92.5005
R512 VDD.n4929 VDD.n4928 92.5005
R513 VDD.n4934 VDD.n4933 92.5005
R514 VDD.n4954 VDD.n4953 92.5005
R515 VDD.n4977 VDD.n4976 92.5005
R516 VDD.n5001 VDD.n5000 92.5005
R517 VDD.n5022 VDD.n5021 92.5005
R518 VDD.n5041 VDD.n5040 92.5005
R519 VDD.n5061 VDD.n5060 92.5005
R520 VDD.n5081 VDD.n5080 92.5005
R521 VDD.n6471 VDD.n6470 92.5005
R522 VDD.n6475 VDD.n6474 92.5005
R523 VDD.n6479 VDD.n6478 92.5005
R524 VDD.n6483 VDD.n6482 92.5005
R525 VDD.n2783 VDD.n2782 92.5005
R526 VDD.n2828 VDD.n2827 92.5005
R527 VDD.n1058 VDD.n1057 92.5005
R528 VDD.n1062 VDD.n1061 92.5005
R529 VDD.n1066 VDD.n1065 92.5005
R530 VDD.n1070 VDD.n1069 92.5005
R531 VDD.n1074 VDD.n1073 92.5005
R532 VDD.n1078 VDD.n1077 92.5005
R533 VDD.n3522 VDD.n3521 92.5005
R534 VDD.n3530 VDD.n3529 92.5005
R535 VDD.n3882 VDD.n3881 92.5005
R536 VDD.n3892 VDD.n3891 92.5005
R537 VDD.n4225 VDD.n4224 92.5005
R538 VDD.n4227 VDD.n4226 92.5005
R539 VDD.n4553 VDD.n4552 92.5005
R540 VDD.n4555 VDD.n4554 92.5005
R541 VDD.n4908 VDD.n4907 92.5005
R542 VDD.n4910 VDD.n4909 92.5005
R543 VDD.n1519 VDD.n1516 92.5005
R544 VDD.n87 VDD.n86 92.5005
R545 VDD.n89 VDD.n88 92.5005
R546 VDD.n9 VDD.n8 92.5005
R547 VDD.n7 VDD.n6 92.5005
R548 VDD.n5 VDD.n4 92.5005
R549 VDD.n3 VDD.n2 92.5005
R550 VDD.n1 VDD.n0 92.5005
R551 VDD.n1518 VDD.n1517 92.5005
R552 VDD.n1565 VDD.n1564 92.5005
R553 VDD.n1563 VDD.n1562 92.5005
R554 VDD.n1560 VDD.n1559 92.5005
R555 VDD.n1558 VDD.n1557 92.5005
R556 VDD.n1556 VDD.n1555 92.5005
R557 VDD.n1571 VDD.n1570 92.5005
R558 VDD.n1547 VDD.n1546 92.5005
R559 VDD.n1545 VDD.n1544 92.5005
R560 VDD.n1542 VDD.n1541 92.5005
R561 VDD.n1540 VDD.n1539 92.5005
R562 VDD.n1538 VDD.n1537 92.5005
R563 VDD.n1553 VDD.n1552 92.5005
R564 VDD.n1681 VDD.n1680 92.5005
R565 VDD.n1679 VDD.n1678 92.5005
R566 VDD.n1676 VDD.n1675 92.5005
R567 VDD.n1674 VDD.n1673 92.5005
R568 VDD.n1672 VDD.n1671 92.5005
R569 VDD.n1687 VDD.n1686 92.5005
R570 VDD.n1703 VDD.n1702 92.5005
R571 VDD.n1701 VDD.n1700 92.5005
R572 VDD.n1698 VDD.n1697 92.5005
R573 VDD.n1696 VDD.n1695 92.5005
R574 VDD.n1694 VDD.n1693 92.5005
R575 VDD.n1709 VDD.n1708 92.5005
R576 VDD.n1246 VDD.n1245 92.5005
R577 VDD.n1244 VDD.n1243 92.5005
R578 VDD.n1241 VDD.n1240 92.5005
R579 VDD.n1239 VDD.n1238 92.5005
R580 VDD.n1237 VDD.n1236 92.5005
R581 VDD.n1252 VDD.n1251 92.5005
R582 VDD.n1234 VDD.n1233 92.5005
R583 VDD.n1228 VDD.n1227 92.5005
R584 VDD.n1226 VDD.n1225 92.5005
R585 VDD.n1223 VDD.n1222 92.5005
R586 VDD.n1322 VDD.n1321 92.5005
R587 VDD.n1325 VDD.n1324 92.5005
R588 VDD.n1428 VDD.n1427 92.5005
R589 VDD.n1424 VDD.n1423 92.5005
R590 VDD.n1422 VDD.n1421 92.5005
R591 VDD.n1419 VDD.n1418 92.5005
R592 VDD.n1417 VDD.n1416 92.5005
R593 VDD.n1414 VDD.n1413 92.5005
R594 VDD.n1381 VDD.n1380 92.5005
R595 VDD.n1430 VDD.n1429 92.5005
R596 VDD.n1433 VDD.n1432 92.5005
R597 VDD.n1436 VDD.n1435 92.5005
R598 VDD.n1439 VDD.n1438 92.5005
R599 VDD.n1445 VDD.n1444 92.5005
R600 VDD.n1412 VDD.n1411 92.5005
R601 VDD.n1410 VDD.n1409 92.5005
R602 VDD.n1408 VDD.n1407 92.5005
R603 VDD.n1406 VDD.n1405 92.5005
R604 VDD.n1404 VDD.n1403 92.5005
R605 VDD.n1402 VDD.n1401 92.5005
R606 VDD.n1399 VDD.n1398 92.5005
R607 VDD.n1397 VDD.n1396 92.5005
R608 VDD.n1395 VDD.n1394 92.5005
R609 VDD.n1393 VDD.n1392 92.5005
R610 VDD.n1391 VDD.n1390 92.5005
R611 VDD.n1389 VDD.n1388 92.5005
R612 VDD.n1386 VDD.n1385 92.5005
R613 VDD.n1590 VDD.n1589 92.5005
R614 VDD.n1596 VDD.n1595 92.5005
R615 VDD.n1602 VDD.n1601 92.5005
R616 VDD.n1608 VDD.n1607 92.5005
R617 VDD.n1614 VDD.n1613 92.5005
R618 VDD.n1627 VDD.n1626 92.5005
R619 VDD.n1633 VDD.n1632 92.5005
R620 VDD.n1639 VDD.n1638 92.5005
R621 VDD.n1645 VDD.n1644 92.5005
R622 VDD.n1651 VDD.n1650 92.5005
R623 VDD.n1657 VDD.n1656 92.5005
R624 VDD.n1783 VDD.n1782 92.5005
R625 VDD.n1777 VDD.n1776 92.5005
R626 VDD.n1771 VDD.n1770 92.5005
R627 VDD.n1765 VDD.n1764 92.5005
R628 VDD.n1759 VDD.n1758 92.5005
R629 VDD.n1753 VDD.n1752 92.5005
R630 VDD.n1740 VDD.n1739 92.5005
R631 VDD.n1734 VDD.n1733 92.5005
R632 VDD.n1728 VDD.n1727 92.5005
R633 VDD.n1329 VDD.n1328 92.5005
R634 VDD.n1331 VDD.n1330 92.5005
R635 VDD.n1333 VDD.n1332 92.5005
R636 VDD.n1336 VDD.n1335 92.5005
R637 VDD.n1338 VDD.n1337 92.5005
R638 VDD.n1340 VDD.n1339 92.5005
R639 VDD.n1342 VDD.n1341 92.5005
R640 VDD.n1344 VDD.n1343 92.5005
R641 VDD.n1346 VDD.n1345 92.5005
R642 VDD.n1349 VDD.n1348 92.5005
R643 VDD.n1351 VDD.n1350 92.5005
R644 VDD.n1353 VDD.n1352 92.5005
R645 VDD.n1355 VDD.n1354 92.5005
R646 VDD.n1371 VDD.n1370 92.5005
R647 VDD.n1367 VDD.n1366 92.5005
R648 VDD.n1365 VDD.n1364 92.5005
R649 VDD.n1362 VDD.n1361 92.5005
R650 VDD.n1360 VDD.n1359 92.5005
R651 VDD.n1357 VDD.n1356 92.5005
R652 VDD.n1505 VDD.n1504 92.5005
R653 VDD.n1504 VDD.n1503 92.5005
R654 VDD.n1500 VDD.n1499 92.5005
R655 VDD.n1499 VDD.n1498 92.5005
R656 VDD.n1495 VDD.n1494 92.5005
R657 VDD.n1494 VDD.n1493 92.5005
R658 VDD.n1490 VDD.n1489 92.5005
R659 VDD.n1489 VDD.n1488 92.5005
R660 VDD.n1485 VDD.n1484 92.5005
R661 VDD.n1484 VDD.n1483 92.5005
R662 VDD.n1480 VDD.n1479 92.5005
R663 VDD.n1479 VDD.n1478 92.5005
R664 VDD.n1470 VDD.n1469 92.5005
R665 VDD.n1469 VDD.n1468 92.5005
R666 VDD.n1465 VDD.n1464 92.5005
R667 VDD.n1464 VDD.n1463 92.5005
R668 VDD.n1460 VDD.n1459 92.5005
R669 VDD.n1459 VDD.n1458 92.5005
R670 VDD.n1455 VDD.n1454 92.5005
R671 VDD.n1454 VDD.n1453 92.5005
R672 VDD.n1450 VDD.n1449 92.5005
R673 VDD.n1449 VDD.n1448 92.5005
R674 VDD.n1574 VDD.n1573 92.5005
R675 VDD.n1573 VDD.n1572 92.5005
R676 VDD.n1586 VDD.n1585 92.5005
R677 VDD.n1585 VDD.n1584 92.5005
R678 VDD.n1592 VDD.n1591 92.5005
R679 VDD.n1591 VDD.n1590 92.5005
R680 VDD.n1598 VDD.n1597 92.5005
R681 VDD.n1597 VDD.n1596 92.5005
R682 VDD.n1604 VDD.n1603 92.5005
R683 VDD.n1603 VDD.n1602 92.5005
R684 VDD.n1610 VDD.n1609 92.5005
R685 VDD.n1609 VDD.n1608 92.5005
R686 VDD.n1616 VDD.n1615 92.5005
R687 VDD.n1615 VDD.n1614 92.5005
R688 VDD.n1629 VDD.n1628 92.5005
R689 VDD.n1628 VDD.n1627 92.5005
R690 VDD.n1635 VDD.n1634 92.5005
R691 VDD.n1634 VDD.n1633 92.5005
R692 VDD.n1641 VDD.n1640 92.5005
R693 VDD.n1640 VDD.n1639 92.5005
R694 VDD.n1647 VDD.n1646 92.5005
R695 VDD.n1646 VDD.n1645 92.5005
R696 VDD.n1653 VDD.n1652 92.5005
R697 VDD.n1652 VDD.n1651 92.5005
R698 VDD.n1659 VDD.n1658 92.5005
R699 VDD.n1658 VDD.n1657 92.5005
R700 VDD.n1785 VDD.n1784 92.5005
R701 VDD.n1784 VDD.n1783 92.5005
R702 VDD.n1779 VDD.n1778 92.5005
R703 VDD.n1778 VDD.n1777 92.5005
R704 VDD.n1773 VDD.n1772 92.5005
R705 VDD.n1772 VDD.n1771 92.5005
R706 VDD.n1767 VDD.n1766 92.5005
R707 VDD.n1766 VDD.n1765 92.5005
R708 VDD.n1761 VDD.n1760 92.5005
R709 VDD.n1760 VDD.n1759 92.5005
R710 VDD.n1755 VDD.n1754 92.5005
R711 VDD.n1754 VDD.n1753 92.5005
R712 VDD.n1742 VDD.n1741 92.5005
R713 VDD.n1741 VDD.n1740 92.5005
R714 VDD.n1736 VDD.n1735 92.5005
R715 VDD.n1735 VDD.n1734 92.5005
R716 VDD.n1730 VDD.n1729 92.5005
R717 VDD.n1729 VDD.n1728 92.5005
R718 VDD.n1724 VDD.n1723 92.5005
R719 VDD.n1723 VDD.n1722 92.5005
R720 VDD.n1719 VDD.n1718 92.5005
R721 VDD.n1718 VDD.n1717 92.5005
R722 VDD.n1714 VDD.n1713 92.5005
R723 VDD.n1713 VDD.n1712 92.5005
R724 VDD.n1260 VDD.n1259 92.5005
R725 VDD.n1259 VDD.n1258 92.5005
R726 VDD.n1265 VDD.n1264 92.5005
R727 VDD.n1264 VDD.n1263 92.5005
R728 VDD.n1270 VDD.n1269 92.5005
R729 VDD.n1269 VDD.n1268 92.5005
R730 VDD.n1275 VDD.n1274 92.5005
R731 VDD.n1274 VDD.n1273 92.5005
R732 VDD.n1280 VDD.n1279 92.5005
R733 VDD.n1279 VDD.n1278 92.5005
R734 VDD.n1285 VDD.n1284 92.5005
R735 VDD.n1284 VDD.n1283 92.5005
R736 VDD.n1312 VDD.n1311 92.5005
R737 VDD.n1311 VDD.n1310 92.5005
R738 VDD.n1307 VDD.n1306 92.5005
R739 VDD.n1306 VDD.n1305 92.5005
R740 VDD.n1302 VDD.n1301 92.5005
R741 VDD.n1301 VDD.n1300 92.5005
R742 VDD.n1297 VDD.n1296 92.5005
R743 VDD.n1296 VDD.n1295 92.5005
R744 VDD.n1082 VDD.n1081 92.5005
R745 VDD.n1091 VDD.n1090 92.5005
R746 VDD.n1093 VDD.n1092 92.5005
R747 VDD.n1087 VDD.n1086 92.5005
R748 VDD.n1521 VDD.n1520 92.5005
R749 VDD.n1523 VDD.n1522 92.5005
R750 VDD.n1514 VDD.n1513 92.5005
R751 VDD.n1512 VDD.n1511 92.5005
R752 VDD.n1509 VDD.n1508 92.5005
R753 VDD.n1507 VDD.n1506 92.5005
R754 VDD.n1502 VDD.n1501 92.5005
R755 VDD.n1497 VDD.n1496 92.5005
R756 VDD.n1492 VDD.n1491 92.5005
R757 VDD.n1487 VDD.n1486 92.5005
R758 VDD.n1482 VDD.n1481 92.5005
R759 VDD.n1477 VDD.n1476 92.5005
R760 VDD.n1475 VDD.n1474 92.5005
R761 VDD.n1472 VDD.n1471 92.5005
R762 VDD.n1467 VDD.n1466 92.5005
R763 VDD.n1462 VDD.n1461 92.5005
R764 VDD.n1457 VDD.n1456 92.5005
R765 VDD.n1452 VDD.n1451 92.5005
R766 VDD.n1447 VDD.n1446 92.5005
R767 VDD.n1576 VDD.n1575 92.5005
R768 VDD.n1578 VDD.n1577 92.5005
R769 VDD.n1581 VDD.n1580 92.5005
R770 VDD.n1583 VDD.n1582 92.5005
R771 VDD.n1588 VDD.n1587 92.5005
R772 VDD.n1594 VDD.n1593 92.5005
R773 VDD.n1600 VDD.n1599 92.5005
R774 VDD.n1606 VDD.n1605 92.5005
R775 VDD.n1612 VDD.n1611 92.5005
R776 VDD.n1618 VDD.n1617 92.5005
R777 VDD.n1620 VDD.n1619 92.5005
R778 VDD.n1623 VDD.n1622 92.5005
R779 VDD.n1625 VDD.n1624 92.5005
R780 VDD.n1631 VDD.n1630 92.5005
R781 VDD.n1637 VDD.n1636 92.5005
R782 VDD.n1643 VDD.n1642 92.5005
R783 VDD.n1649 VDD.n1648 92.5005
R784 VDD.n1655 VDD.n1654 92.5005
R785 VDD.n1792 VDD.n1791 92.5005
R786 VDD.n1789 VDD.n1788 92.5005
R787 VDD.n1787 VDD.n1786 92.5005
R788 VDD.n1781 VDD.n1780 92.5005
R789 VDD.n1775 VDD.n1774 92.5005
R790 VDD.n1769 VDD.n1768 92.5005
R791 VDD.n1763 VDD.n1762 92.5005
R792 VDD.n1757 VDD.n1756 92.5005
R793 VDD.n1751 VDD.n1750 92.5005
R794 VDD.n1749 VDD.n1748 92.5005
R795 VDD.n1746 VDD.n1745 92.5005
R796 VDD.n1744 VDD.n1743 92.5005
R797 VDD.n1738 VDD.n1737 92.5005
R798 VDD.n1732 VDD.n1731 92.5005
R799 VDD.n1726 VDD.n1725 92.5005
R800 VDD.n1721 VDD.n1720 92.5005
R801 VDD.n1716 VDD.n1715 92.5005
R802 VDD.n1711 VDD.n1710 92.5005
R803 VDD.n1254 VDD.n1253 92.5005
R804 VDD.n1257 VDD.n1256 92.5005
R805 VDD.n1262 VDD.n1261 92.5005
R806 VDD.n1267 VDD.n1266 92.5005
R807 VDD.n1272 VDD.n1271 92.5005
R808 VDD.n1277 VDD.n1276 92.5005
R809 VDD.n1282 VDD.n1281 92.5005
R810 VDD.n1287 VDD.n1286 92.5005
R811 VDD.n1289 VDD.n1288 92.5005
R812 VDD.n1292 VDD.n1291 92.5005
R813 VDD.n1294 VDD.n1293 92.5005
R814 VDD.n1299 VDD.n1298 92.5005
R815 VDD.n1304 VDD.n1303 92.5005
R816 VDD.n1309 VDD.n1308 92.5005
R817 VDD.n1314 VDD.n1313 92.5005
R818 VDD.n1317 VDD.n1316 92.5005
R819 VDD.n1319 VDD.n1318 92.5005
R820 VDD.n1221 VDD.n1220 92.5005
R821 VDD.n1219 VDD.n1218 92.5005
R822 VDD.n1217 VDD.n1216 92.5005
R823 VDD.n1215 VDD.n1214 92.5005
R824 VDD.n1213 VDD.n1212 92.5005
R825 VDD.n1211 VDD.n1210 92.5005
R826 VDD.n1195 VDD.n1194 92.5005
R827 VDD.n1197 VDD.n1196 92.5005
R828 VDD.n1199 VDD.n1198 92.5005
R829 VDD.n1201 VDD.n1200 92.5005
R830 VDD.n1203 VDD.n1202 92.5005
R831 VDD.n1205 VDD.n1204 92.5005
R832 VDD.n1193 VDD.n1192 92.5005
R833 VDD.n1191 VDD.n1190 92.5005
R834 VDD.n1103 VDD.n1095 92.5005
R835 VDD.n1097 VDD.n1096 92.5005
R836 VDD.n1099 VDD.n1098 92.5005
R837 VDD.n1084 VDD.n1083 92.5005
R838 VDD.n1103 VDD.n1102 92.5005
R839 VDD.n1102 VDD.n1101 92.5005
R840 VDD.n1158 VDD.n1157 92.5005
R841 VDD.n1157 VDD.n1156 92.5005
R842 VDD.n1161 VDD.n1160 92.5005
R843 VDD.n1160 VDD.n1159 92.5005
R844 VDD.n1164 VDD.n1163 92.5005
R845 VDD.n1163 VDD.n1162 92.5005
R846 VDD.n1167 VDD.n1166 92.5005
R847 VDD.n1166 VDD.n1165 92.5005
R848 VDD.n1170 VDD.n1169 92.5005
R849 VDD.n1169 VDD.n1168 92.5005
R850 VDD.n1173 VDD.n1172 92.5005
R851 VDD.n1172 VDD.n1171 92.5005
R852 VDD.n1176 VDD.n1175 92.5005
R853 VDD.n1175 VDD.n1174 92.5005
R854 VDD.n1179 VDD.n1178 92.5005
R855 VDD.n1178 VDD.n1177 92.5005
R856 VDD.n1182 VDD.n1181 92.5005
R857 VDD.n1181 VDD.n1180 92.5005
R858 VDD.n1185 VDD.n1184 92.5005
R859 VDD.n1184 VDD.n1183 92.5005
R860 VDD.n1188 VDD.n1187 92.5005
R861 VDD.n1187 VDD.n1186 92.5005
R862 VDD.n868 VDD.n867 92.5005
R863 VDD.n161 VDD.n160 92.5005
R864 VDD.n882 VDD.n881 92.5005
R865 VDD.n885 VDD.n884 92.5005
R866 VDD.n884 VDD.n883 92.5005
R867 VDD.n889 VDD.n888 92.5005
R868 VDD.n888 VDD.n887 92.5005
R869 VDD.n119 VDD.n118 92.5005
R870 VDD.n118 VDD.n117 92.5005
R871 VDD.n131 VDD.n130 92.5005
R872 VDD.n130 VDD.n129 92.5005
R873 VDD.n899 VDD.n898 92.5005
R874 VDD.n898 VDD.n897 92.5005
R875 VDD.n895 VDD.n894 92.5005
R876 VDD.n894 VDD.n893 92.5005
R877 VDD.n907 VDD.n906 92.5005
R878 VDD.n906 VDD.n905 92.5005
R879 VDD.n912 VDD.n911 92.5005
R880 VDD.n911 VDD.n910 92.5005
R881 VDD.n920 VDD.n919 92.5005
R882 VDD.n919 VDD.n918 92.5005
R883 VDD.n917 VDD.n916 92.5005
R884 VDD.n916 VDD.n915 92.5005
R885 VDD.n925 VDD.n924 92.5005
R886 VDD.n924 VDD.n923 92.5005
R887 VDD.n930 VDD.n929 92.5005
R888 VDD.n929 VDD.n928 92.5005
R889 VDD.n935 VDD.n934 92.5005
R890 VDD.n934 VDD.n933 92.5005
R891 VDD.n940 VDD.n939 92.5005
R892 VDD.n939 VDD.n938 92.5005
R893 VDD.n945 VDD.n944 92.5005
R894 VDD.n944 VDD.n943 92.5005
R895 VDD.n1016 VDD.n1015 92.5005
R896 VDD.n1015 VDD.n1014 92.5005
R897 VDD.n1013 VDD.n1012 92.5005
R898 VDD.n1012 VDD.n1011 92.5005
R899 VDD.n1010 VDD.n1009 92.5005
R900 VDD.n1009 VDD.n1008 92.5005
R901 VDD.n1007 VDD.n1006 92.5005
R902 VDD.n1006 VDD.n1005 92.5005
R903 VDD.n1004 VDD.n1003 92.5005
R904 VDD.n1003 VDD.n1002 92.5005
R905 VDD.n1001 VDD.n1000 92.5005
R906 VDD.n1000 VDD.n999 92.5005
R907 VDD.n998 VDD.n997 92.5005
R908 VDD.n997 VDD.n996 92.5005
R909 VDD.n995 VDD.n994 92.5005
R910 VDD.n994 VDD.n993 92.5005
R911 VDD.n992 VDD.n991 92.5005
R912 VDD.n991 VDD.n990 92.5005
R913 VDD.n989 VDD.n988 92.5005
R914 VDD.n988 VDD.n987 92.5005
R915 VDD.n986 VDD.n985 92.5005
R916 VDD.n985 VDD.n984 92.5005
R917 VDD.n983 VDD.n982 92.5005
R918 VDD.n982 VDD.n981 92.5005
R919 VDD.n980 VDD.n979 92.5005
R920 VDD.n979 VDD.n978 92.5005
R921 VDD.n977 VDD.n976 92.5005
R922 VDD.n976 VDD.n975 92.5005
R923 VDD.n974 VDD.n973 92.5005
R924 VDD.n973 VDD.n972 92.5005
R925 VDD.n971 VDD.n970 92.5005
R926 VDD.n970 VDD.n969 92.5005
R927 VDD.n968 VDD.n967 92.5005
R928 VDD.n967 VDD.n966 92.5005
R929 VDD.n965 VDD.n964 92.5005
R930 VDD.n964 VDD.n963 92.5005
R931 VDD.n962 VDD.n961 92.5005
R932 VDD.n961 VDD.n960 92.5005
R933 VDD.n959 VDD.n958 92.5005
R934 VDD.n958 VDD.n957 92.5005
R935 VDD.n956 VDD.n955 92.5005
R936 VDD.n955 VDD.n954 92.5005
R937 VDD.n953 VDD.n952 92.5005
R938 VDD.n952 VDD.n951 92.5005
R939 VDD.n950 VDD.n949 92.5005
R940 VDD.n949 VDD.n948 92.5005
R941 VDD.n1107 VDD.n1106 92.5005
R942 VDD.n1106 VDD.n1105 92.5005
R943 VDD.n1110 VDD.n1109 92.5005
R944 VDD.n1109 VDD.n1108 92.5005
R945 VDD.n1113 VDD.n1112 92.5005
R946 VDD.n1112 VDD.n1111 92.5005
R947 VDD.n1116 VDD.n1115 92.5005
R948 VDD.n1115 VDD.n1114 92.5005
R949 VDD.n1119 VDD.n1118 92.5005
R950 VDD.n1118 VDD.n1117 92.5005
R951 VDD.n1122 VDD.n1121 92.5005
R952 VDD.n1121 VDD.n1120 92.5005
R953 VDD.n1125 VDD.n1124 92.5005
R954 VDD.n1124 VDD.n1123 92.5005
R955 VDD.n1128 VDD.n1127 92.5005
R956 VDD.n1127 VDD.n1126 92.5005
R957 VDD.n1131 VDD.n1130 92.5005
R958 VDD.n1130 VDD.n1129 92.5005
R959 VDD.n1134 VDD.n1133 92.5005
R960 VDD.n1133 VDD.n1132 92.5005
R961 VDD.n1137 VDD.n1136 92.5005
R962 VDD.n1136 VDD.n1135 92.5005
R963 VDD.n1140 VDD.n1139 92.5005
R964 VDD.n1139 VDD.n1138 92.5005
R965 VDD.n1143 VDD.n1142 92.5005
R966 VDD.n1142 VDD.n1141 92.5005
R967 VDD.n1146 VDD.n1145 92.5005
R968 VDD.n1145 VDD.n1144 92.5005
R969 VDD.n1149 VDD.n1148 92.5005
R970 VDD.n1148 VDD.n1147 92.5005
R971 VDD.n1152 VDD.n1151 92.5005
R972 VDD.n1151 VDD.n1150 92.5005
R973 VDD.n1155 VDD.n1154 92.5005
R974 VDD.n1154 VDD.n1153 92.5005
R975 VDD.n870 VDD.n869 92.5005
R976 VDD.n873 VDD.n872 92.5005
R977 VDD.n379 VDD.n378 92.5005
R978 VDD.n378 VDD.n377 92.5005
R979 VDD.n384 VDD.n383 92.5005
R980 VDD.n383 VDD.n382 92.5005
R981 VDD.n389 VDD.n388 92.5005
R982 VDD.n388 VDD.n387 92.5005
R983 VDD.n397 VDD.n396 92.5005
R984 VDD.n396 VDD.n395 92.5005
R985 VDD.n394 VDD.n393 92.5005
R986 VDD.n393 VDD.n392 92.5005
R987 VDD.n402 VDD.n401 92.5005
R988 VDD.n401 VDD.n400 92.5005
R989 VDD.n407 VDD.n406 92.5005
R990 VDD.n406 VDD.n405 92.5005
R991 VDD.n412 VDD.n411 92.5005
R992 VDD.n411 VDD.n410 92.5005
R993 VDD.n417 VDD.n416 92.5005
R994 VDD.n416 VDD.n415 92.5005
R995 VDD.n422 VDD.n421 92.5005
R996 VDD.n421 VDD.n420 92.5005
R997 VDD.n427 VDD.n426 92.5005
R998 VDD.n426 VDD.n425 92.5005
R999 VDD.n432 VDD.n431 92.5005
R1000 VDD.n431 VDD.n430 92.5005
R1001 VDD.n437 VDD.n436 92.5005
R1002 VDD.n436 VDD.n435 92.5005
R1003 VDD.n442 VDD.n441 92.5005
R1004 VDD.n441 VDD.n440 92.5005
R1005 VDD.n447 VDD.n446 92.5005
R1006 VDD.n446 VDD.n445 92.5005
R1007 VDD.n452 VDD.n451 92.5005
R1008 VDD.n451 VDD.n450 92.5005
R1009 VDD.n457 VDD.n456 92.5005
R1010 VDD.n456 VDD.n455 92.5005
R1011 VDD.n462 VDD.n461 92.5005
R1012 VDD.n461 VDD.n460 92.5005
R1013 VDD.n467 VDD.n466 92.5005
R1014 VDD.n466 VDD.n465 92.5005
R1015 VDD.n472 VDD.n471 92.5005
R1016 VDD.n471 VDD.n470 92.5005
R1017 VDD.n477 VDD.n476 92.5005
R1018 VDD.n476 VDD.n475 92.5005
R1019 VDD.n485 VDD.n484 92.5005
R1020 VDD.n484 VDD.n483 92.5005
R1021 VDD.n482 VDD.n481 92.5005
R1022 VDD.n481 VDD.n480 92.5005
R1023 VDD.n490 VDD.n489 92.5005
R1024 VDD.n489 VDD.n488 92.5005
R1025 VDD.n495 VDD.n494 92.5005
R1026 VDD.n494 VDD.n493 92.5005
R1027 VDD.n500 VDD.n499 92.5005
R1028 VDD.n499 VDD.n498 92.5005
R1029 VDD.n505 VDD.n504 92.5005
R1030 VDD.n504 VDD.n503 92.5005
R1031 VDD.n510 VDD.n509 92.5005
R1032 VDD.n509 VDD.n508 92.5005
R1033 VDD.n515 VDD.n514 92.5005
R1034 VDD.n514 VDD.n513 92.5005
R1035 VDD.n520 VDD.n519 92.5005
R1036 VDD.n519 VDD.n518 92.5005
R1037 VDD.n525 VDD.n524 92.5005
R1038 VDD.n524 VDD.n523 92.5005
R1039 VDD.n530 VDD.n529 92.5005
R1040 VDD.n529 VDD.n528 92.5005
R1041 VDD.n535 VDD.n534 92.5005
R1042 VDD.n534 VDD.n533 92.5005
R1043 VDD.n540 VDD.n539 92.5005
R1044 VDD.n539 VDD.n538 92.5005
R1045 VDD.n545 VDD.n544 92.5005
R1046 VDD.n544 VDD.n543 92.5005
R1047 VDD.n550 VDD.n549 92.5005
R1048 VDD.n549 VDD.n548 92.5005
R1049 VDD.n555 VDD.n554 92.5005
R1050 VDD.n554 VDD.n553 92.5005
R1051 VDD.n560 VDD.n559 92.5005
R1052 VDD.n559 VDD.n558 92.5005
R1053 VDD.n565 VDD.n564 92.5005
R1054 VDD.n564 VDD.n563 92.5005
R1055 VDD.n573 VDD.n572 92.5005
R1056 VDD.n572 VDD.n571 92.5005
R1057 VDD.n570 VDD.n569 92.5005
R1058 VDD.n569 VDD.n568 92.5005
R1059 VDD.n578 VDD.n577 92.5005
R1060 VDD.n577 VDD.n576 92.5005
R1061 VDD.n583 VDD.n582 92.5005
R1062 VDD.n582 VDD.n581 92.5005
R1063 VDD.n588 VDD.n587 92.5005
R1064 VDD.n587 VDD.n586 92.5005
R1065 VDD.n593 VDD.n592 92.5005
R1066 VDD.n592 VDD.n591 92.5005
R1067 VDD.n598 VDD.n597 92.5005
R1068 VDD.n597 VDD.n596 92.5005
R1069 VDD.n603 VDD.n602 92.5005
R1070 VDD.n602 VDD.n601 92.5005
R1071 VDD.n608 VDD.n607 92.5005
R1072 VDD.n607 VDD.n606 92.5005
R1073 VDD.n613 VDD.n612 92.5005
R1074 VDD.n612 VDD.n611 92.5005
R1075 VDD.n618 VDD.n617 92.5005
R1076 VDD.n617 VDD.n616 92.5005
R1077 VDD.n623 VDD.n622 92.5005
R1078 VDD.n622 VDD.n621 92.5005
R1079 VDD.n628 VDD.n627 92.5005
R1080 VDD.n627 VDD.n626 92.5005
R1081 VDD.n633 VDD.n632 92.5005
R1082 VDD.n632 VDD.n631 92.5005
R1083 VDD.n638 VDD.n637 92.5005
R1084 VDD.n637 VDD.n636 92.5005
R1085 VDD.n643 VDD.n642 92.5005
R1086 VDD.n642 VDD.n641 92.5005
R1087 VDD.n648 VDD.n647 92.5005
R1088 VDD.n647 VDD.n646 92.5005
R1089 VDD.n653 VDD.n652 92.5005
R1090 VDD.n652 VDD.n651 92.5005
R1091 VDD.n661 VDD.n660 92.5005
R1092 VDD.n660 VDD.n659 92.5005
R1093 VDD.n658 VDD.n657 92.5005
R1094 VDD.n657 VDD.n656 92.5005
R1095 VDD.n666 VDD.n665 92.5005
R1096 VDD.n665 VDD.n664 92.5005
R1097 VDD.n671 VDD.n670 92.5005
R1098 VDD.n670 VDD.n669 92.5005
R1099 VDD.n676 VDD.n675 92.5005
R1100 VDD.n675 VDD.n674 92.5005
R1101 VDD.n681 VDD.n680 92.5005
R1102 VDD.n680 VDD.n679 92.5005
R1103 VDD.n686 VDD.n685 92.5005
R1104 VDD.n685 VDD.n684 92.5005
R1105 VDD.n691 VDD.n690 92.5005
R1106 VDD.n690 VDD.n689 92.5005
R1107 VDD.n696 VDD.n695 92.5005
R1108 VDD.n695 VDD.n694 92.5005
R1109 VDD.n701 VDD.n700 92.5005
R1110 VDD.n700 VDD.n699 92.5005
R1111 VDD.n706 VDD.n705 92.5005
R1112 VDD.n705 VDD.n704 92.5005
R1113 VDD.n711 VDD.n710 92.5005
R1114 VDD.n710 VDD.n709 92.5005
R1115 VDD.n716 VDD.n715 92.5005
R1116 VDD.n715 VDD.n714 92.5005
R1117 VDD.n721 VDD.n720 92.5005
R1118 VDD.n720 VDD.n719 92.5005
R1119 VDD.n726 VDD.n725 92.5005
R1120 VDD.n725 VDD.n724 92.5005
R1121 VDD.n731 VDD.n730 92.5005
R1122 VDD.n730 VDD.n729 92.5005
R1123 VDD.n736 VDD.n735 92.5005
R1124 VDD.n735 VDD.n734 92.5005
R1125 VDD.n741 VDD.n740 92.5005
R1126 VDD.n740 VDD.n739 92.5005
R1127 VDD.n749 VDD.n748 92.5005
R1128 VDD.n748 VDD.n747 92.5005
R1129 VDD.n746 VDD.n745 92.5005
R1130 VDD.n745 VDD.n744 92.5005
R1131 VDD.n754 VDD.n753 92.5005
R1132 VDD.n753 VDD.n752 92.5005
R1133 VDD.n759 VDD.n758 92.5005
R1134 VDD.n758 VDD.n757 92.5005
R1135 VDD.n764 VDD.n763 92.5005
R1136 VDD.n763 VDD.n762 92.5005
R1137 VDD.n769 VDD.n768 92.5005
R1138 VDD.n768 VDD.n767 92.5005
R1139 VDD.n774 VDD.n773 92.5005
R1140 VDD.n773 VDD.n772 92.5005
R1141 VDD.n779 VDD.n778 92.5005
R1142 VDD.n778 VDD.n777 92.5005
R1143 VDD.n784 VDD.n783 92.5005
R1144 VDD.n783 VDD.n782 92.5005
R1145 VDD.n789 VDD.n788 92.5005
R1146 VDD.n788 VDD.n787 92.5005
R1147 VDD.n794 VDD.n793 92.5005
R1148 VDD.n793 VDD.n792 92.5005
R1149 VDD.n799 VDD.n798 92.5005
R1150 VDD.n798 VDD.n797 92.5005
R1151 VDD.n804 VDD.n803 92.5005
R1152 VDD.n803 VDD.n802 92.5005
R1153 VDD.n809 VDD.n808 92.5005
R1154 VDD.n808 VDD.n807 92.5005
R1155 VDD.n814 VDD.n813 92.5005
R1156 VDD.n813 VDD.n812 92.5005
R1157 VDD.n819 VDD.n818 92.5005
R1158 VDD.n818 VDD.n817 92.5005
R1159 VDD.n824 VDD.n823 92.5005
R1160 VDD.n823 VDD.n822 92.5005
R1161 VDD.n829 VDD.n828 92.5005
R1162 VDD.n828 VDD.n827 92.5005
R1163 VDD.n837 VDD.n836 92.5005
R1164 VDD.n836 VDD.n835 92.5005
R1165 VDD.n834 VDD.n833 92.5005
R1166 VDD.n833 VDD.n832 92.5005
R1167 VDD.n842 VDD.n841 92.5005
R1168 VDD.n841 VDD.n840 92.5005
R1169 VDD.n847 VDD.n846 92.5005
R1170 VDD.n846 VDD.n845 92.5005
R1171 VDD.n852 VDD.n851 92.5005
R1172 VDD.n851 VDD.n850 92.5005
R1173 VDD.n857 VDD.n856 92.5005
R1174 VDD.n856 VDD.n855 92.5005
R1175 VDD.n862 VDD.n861 92.5005
R1176 VDD.n861 VDD.n860 92.5005
R1177 VDD.n363 VDD.n362 92.5005
R1178 VDD.n6749 VDD.n6748 92.5005
R1179 VDD.n6748 VDD.n6747 92.5005
R1180 VDD.n6746 VDD.n6745 92.5005
R1181 VDD.n6745 VDD.n6744 92.5005
R1182 VDD.n6743 VDD.n6742 92.5005
R1183 VDD.n6742 VDD.n6741 92.5005
R1184 VDD.n6740 VDD.n6739 92.5005
R1185 VDD.n6739 VDD.n6738 92.5005
R1186 VDD.n6737 VDD.n6736 92.5005
R1187 VDD.n6736 VDD.n6735 92.5005
R1188 VDD.n6734 VDD.n6733 92.5005
R1189 VDD.n6733 VDD.n6732 92.5005
R1190 VDD.n6731 VDD.n6730 92.5005
R1191 VDD.n6730 VDD.n6729 92.5005
R1192 VDD.n6728 VDD.n6727 92.5005
R1193 VDD.n6727 VDD.n6726 92.5005
R1194 VDD.n6725 VDD.n6724 92.5005
R1195 VDD.n6724 VDD.n6723 92.5005
R1196 VDD.n6722 VDD.n6721 92.5005
R1197 VDD.n6721 VDD.n6720 92.5005
R1198 VDD.n6719 VDD.n6718 92.5005
R1199 VDD.n6718 VDD.n6717 92.5005
R1200 VDD.n172 VDD.n171 92.5005
R1201 VDD.n171 VDD.n170 92.5005
R1202 VDD.n175 VDD.n174 92.5005
R1203 VDD.n174 VDD.n173 92.5005
R1204 VDD.n179 VDD.n178 92.5005
R1205 VDD.n178 VDD.n177 92.5005
R1206 VDD.n184 VDD.n183 92.5005
R1207 VDD.n183 VDD.n182 92.5005
R1208 VDD.n189 VDD.n188 92.5005
R1209 VDD.n188 VDD.n187 92.5005
R1210 VDD.n194 VDD.n193 92.5005
R1211 VDD.n193 VDD.n192 92.5005
R1212 VDD.n199 VDD.n198 92.5005
R1213 VDD.n198 VDD.n197 92.5005
R1214 VDD.n202 VDD.n201 92.5005
R1215 VDD.n201 VDD.n200 92.5005
R1216 VDD.n207 VDD.n206 92.5005
R1217 VDD.n206 VDD.n205 92.5005
R1218 VDD.n212 VDD.n211 92.5005
R1219 VDD.n211 VDD.n210 92.5005
R1220 VDD.n217 VDD.n216 92.5005
R1221 VDD.n216 VDD.n215 92.5005
R1222 VDD.n222 VDD.n221 92.5005
R1223 VDD.n221 VDD.n220 92.5005
R1224 VDD.n227 VDD.n226 92.5005
R1225 VDD.n226 VDD.n225 92.5005
R1226 VDD.n232 VDD.n231 92.5005
R1227 VDD.n231 VDD.n230 92.5005
R1228 VDD.n237 VDD.n236 92.5005
R1229 VDD.n236 VDD.n235 92.5005
R1230 VDD.n242 VDD.n241 92.5005
R1231 VDD.n241 VDD.n240 92.5005
R1232 VDD.n247 VDD.n246 92.5005
R1233 VDD.n246 VDD.n245 92.5005
R1234 VDD.n252 VDD.n251 92.5005
R1235 VDD.n251 VDD.n250 92.5005
R1236 VDD.n257 VDD.n256 92.5005
R1237 VDD.n256 VDD.n255 92.5005
R1238 VDD.n165 VDD.n164 92.5005
R1239 VDD.n164 VDD.n163 92.5005
R1240 VDD.n169 VDD.n168 92.5005
R1241 VDD.n168 VDD.n167 92.5005
R1242 VDD.n264 VDD.n263 92.5005
R1243 VDD.n263 VDD.n262 92.5005
R1244 VDD.n267 VDD.n266 92.5005
R1245 VDD.n266 VDD.n265 92.5005
R1246 VDD.n270 VDD.n269 92.5005
R1247 VDD.n269 VDD.n268 92.5005
R1248 VDD.n273 VDD.n272 92.5005
R1249 VDD.n272 VDD.n271 92.5005
R1250 VDD.n276 VDD.n275 92.5005
R1251 VDD.n275 VDD.n274 92.5005
R1252 VDD.n279 VDD.n278 92.5005
R1253 VDD.n278 VDD.n277 92.5005
R1254 VDD.n282 VDD.n281 92.5005
R1255 VDD.n281 VDD.n280 92.5005
R1256 VDD.n285 VDD.n284 92.5005
R1257 VDD.n284 VDD.n283 92.5005
R1258 VDD.n288 VDD.n287 92.5005
R1259 VDD.n287 VDD.n286 92.5005
R1260 VDD.n291 VDD.n290 92.5005
R1261 VDD.n290 VDD.n289 92.5005
R1262 VDD.n295 VDD.n294 92.5005
R1263 VDD.n294 VDD.n293 92.5005
R1264 VDD.n300 VDD.n299 92.5005
R1265 VDD.n299 VDD.n298 92.5005
R1266 VDD.n305 VDD.n304 92.5005
R1267 VDD.n304 VDD.n303 92.5005
R1268 VDD.n310 VDD.n309 92.5005
R1269 VDD.n309 VDD.n308 92.5005
R1270 VDD.n315 VDD.n314 92.5005
R1271 VDD.n314 VDD.n313 92.5005
R1272 VDD.n320 VDD.n319 92.5005
R1273 VDD.n319 VDD.n318 92.5005
R1274 VDD.n325 VDD.n324 92.5005
R1275 VDD.n324 VDD.n323 92.5005
R1276 VDD.n330 VDD.n329 92.5005
R1277 VDD.n329 VDD.n328 92.5005
R1278 VDD.n335 VDD.n334 92.5005
R1279 VDD.n334 VDD.n333 92.5005
R1280 VDD.n340 VDD.n339 92.5005
R1281 VDD.n339 VDD.n338 92.5005
R1282 VDD.n343 VDD.n342 92.5005
R1283 VDD.n342 VDD.n341 92.5005
R1284 VDD.n348 VDD.n347 92.5005
R1285 VDD.n347 VDD.n346 92.5005
R1286 VDD.n353 VDD.n352 92.5005
R1287 VDD.n352 VDD.n351 92.5005
R1288 VDD.n359 VDD.n358 92.5005
R1289 VDD.n365 VDD.n364 92.5005
R1290 VDD.n370 VDD.n369 92.5005
R1291 VDD.n372 VDD.n371 92.5005
R1292 VDD.n6786 VDD.n6785 92.5005
R1293 VDD.n6785 VDD.n6784 92.5005
R1294 VDD.n6782 VDD.n6781 92.5005
R1295 VDD.n6781 VDD.n6780 92.5005
R1296 VDD.n6779 VDD.n6778 92.5005
R1297 VDD.n6778 VDD.n6777 92.5005
R1298 VDD.n6776 VDD.n6775 92.5005
R1299 VDD.n6775 VDD.n6774 92.5005
R1300 VDD.n6773 VDD.n6772 92.5005
R1301 VDD.n6772 VDD.n6771 92.5005
R1302 VDD.n6770 VDD.n6769 92.5005
R1303 VDD.n6769 VDD.n6768 92.5005
R1304 VDD.n6767 VDD.n6766 92.5005
R1305 VDD.n6766 VDD.n6765 92.5005
R1306 VDD.n6764 VDD.n6763 92.5005
R1307 VDD.n6763 VDD.n6762 92.5005
R1308 VDD.n6761 VDD.n6760 92.5005
R1309 VDD.n6760 VDD.n6759 92.5005
R1310 VDD.n6758 VDD.n6757 92.5005
R1311 VDD.n6757 VDD.n6756 92.5005
R1312 VDD.n6755 VDD.n6754 92.5005
R1313 VDD.n6754 VDD.n6753 92.5005
R1314 VDD.n6752 VDD.n6751 92.5005
R1315 VDD.n6751 VDD.n6750 92.5005
R1316 VDD.n6789 VDD.n6788 92.5005
R1317 VDD.n6788 VDD.n6787 92.5005
R1318 VDD.n6716 VDD.n6715 92.5005
R1319 VDD.n6715 VDD.n6714 92.5005
R1320 VDD.n6713 VDD.n6712 92.5005
R1321 VDD.n6712 VDD.n6711 92.5005
R1322 VDD.n84 VDD.n83 92.5005
R1323 VDD.n83 VDD.n82 92.5005
R1324 VDD.n81 VDD.n80 92.5005
R1325 VDD.n80 VDD.n79 92.5005
R1326 VDD.n78 VDD.n77 92.5005
R1327 VDD.n77 VDD.n76 92.5005
R1328 VDD.n67 VDD.n66 92.5005
R1329 VDD.n63 VDD.n62 92.5005
R1330 VDD.n59 VDD.n58 92.5005
R1331 VDD.n55 VDD.n54 92.5005
R1332 VDD.n51 VDD.n50 92.5005
R1333 VDD.n47 VDD.n46 92.5005
R1334 VDD.n43 VDD.n42 92.5005
R1335 VDD.n39 VDD.n38 92.5005
R1336 VDD.n35 VDD.n34 92.5005
R1337 VDD.n31 VDD.n30 92.5005
R1338 VDD.n27 VDD.n26 92.5005
R1339 VDD.n23 VDD.n22 92.5005
R1340 VDD.n19 VDD.n18 92.5005
R1341 VDD.n15 VDD.n14 92.5005
R1342 VDD.n11 VDD.n10 92.5005
R1343 VDD.n5284 VDD.n5283 92.5005
R1344 VDD.n5288 VDD.n5287 92.5005
R1345 VDD.n5292 VDD.n5291 92.5005
R1346 VDD.n5296 VDD.n5295 92.5005
R1347 VDD.n5300 VDD.n5299 92.5005
R1348 VDD.n5304 VDD.n5303 92.5005
R1349 VDD.n5308 VDD.n5307 92.5005
R1350 VDD.n5312 VDD.n5311 92.5005
R1351 VDD.n5316 VDD.n5315 92.5005
R1352 VDD.n5320 VDD.n5319 92.5005
R1353 VDD.n5324 VDD.n5323 92.5005
R1354 VDD.n5328 VDD.n5327 92.5005
R1355 VDD.n5332 VDD.n5331 92.5005
R1356 VDD.n5336 VDD.n5335 92.5005
R1357 VDD.n5340 VDD.n5339 92.5005
R1358 VDD.n5344 VDD.n5343 92.5005
R1359 VDD.n5348 VDD.n5347 92.5005
R1360 VDD.n6501 VDD.n6500 92.5005
R1361 VDD.n6503 VDD.n6502 92.5005
R1362 VDD.n6429 VDD.n6428 92.5005
R1363 VDD.n6425 VDD.n6424 92.5005
R1364 VDD.n6419 VDD.n6418 92.5005
R1365 VDD.n6413 VDD.n6412 92.5005
R1366 VDD.n6407 VDD.n6406 92.5005
R1367 VDD.n6401 VDD.n6400 92.5005
R1368 VDD.n6395 VDD.n6394 92.5005
R1369 VDD.n6389 VDD.n6388 92.5005
R1370 VDD.n6383 VDD.n6382 92.5005
R1371 VDD.n6375 VDD.n6374 92.5005
R1372 VDD.n6367 VDD.n6366 92.5005
R1373 VDD.n6359 VDD.n6358 92.5005
R1374 VDD.n6361 VDD.n6360 92.5005
R1375 VDD.n6353 VDD.n6352 92.5005
R1376 VDD.n6347 VDD.n6346 92.5005
R1377 VDD.n6341 VDD.n6340 92.5005
R1378 VDD.n6335 VDD.n6334 92.5005
R1379 VDD.n6329 VDD.n6328 92.5005
R1380 VDD.n6323 VDD.n6322 92.5005
R1381 VDD.n6319 VDD.n6318 92.5005
R1382 VDD.n6313 VDD.n6312 92.5005
R1383 VDD.n6307 VDD.n6306 92.5005
R1384 VDD.n6301 VDD.n6300 92.5005
R1385 VDD.n6295 VDD.n6294 92.5005
R1386 VDD.n6289 VDD.n6288 92.5005
R1387 VDD.n6283 VDD.n6282 92.5005
R1388 VDD.n6277 VDD.n6276 92.5005
R1389 VDD.n6269 VDD.n6268 92.5005
R1390 VDD.n6261 VDD.n6260 92.5005
R1391 VDD.n6271 VDD.n6270 92.5005
R1392 VDD.n6267 VDD.n6266 92.5005
R1393 VDD.n6275 VDD.n6274 92.5005
R1394 VDD.n6281 VDD.n6280 92.5005
R1395 VDD.n6287 VDD.n6286 92.5005
R1396 VDD.n6293 VDD.n6292 92.5005
R1397 VDD.n6299 VDD.n6298 92.5005
R1398 VDD.n6305 VDD.n6304 92.5005
R1399 VDD.n6311 VDD.n6310 92.5005
R1400 VDD.n6317 VDD.n6316 92.5005
R1401 VDD.n6325 VDD.n6324 92.5005
R1402 VDD.n6331 VDD.n6330 92.5005
R1403 VDD.n6337 VDD.n6336 92.5005
R1404 VDD.n6343 VDD.n6342 92.5005
R1405 VDD.n6349 VDD.n6348 92.5005
R1406 VDD.n6355 VDD.n6354 92.5005
R1407 VDD.n6363 VDD.n6362 92.5005
R1408 VDD.n6369 VDD.n6368 92.5005
R1409 VDD.n6377 VDD.n6376 92.5005
R1410 VDD.n6373 VDD.n6372 92.5005
R1411 VDD.n6381 VDD.n6380 92.5005
R1412 VDD.n6387 VDD.n6386 92.5005
R1413 VDD.n6393 VDD.n6392 92.5005
R1414 VDD.n6399 VDD.n6398 92.5005
R1415 VDD.n6405 VDD.n6404 92.5005
R1416 VDD.n6411 VDD.n6410 92.5005
R1417 VDD.n6417 VDD.n6416 92.5005
R1418 VDD.n6423 VDD.n6422 92.5005
R1419 VDD.n6263 VDD.n6262 92.5005
R1420 VDD.n6254 VDD.n6253 92.5005
R1421 VDD.n6258 VDD.n6257 92.5005
R1422 VDD.n6256 VDD.n6255 92.5005
R1423 VDD.n5272 VDD.n5271 92.5005
R1424 VDD.n5274 VDD.n5273 92.5005
R1425 VDD.n5276 VDD.n5275 92.5005
R1426 VDD.n5278 VDD.n5277 92.5005
R1427 VDD.n5280 VDD.n5279 92.5005
R1428 VDD.n5352 VDD.n5351 92.5005
R1429 VDD.n5350 VDD.n5349 92.5005
R1430 VDD.n5346 VDD.n5345 92.5005
R1431 VDD.n5342 VDD.n5341 92.5005
R1432 VDD.n5338 VDD.n5337 92.5005
R1433 VDD.n5334 VDD.n5333 92.5005
R1434 VDD.n5330 VDD.n5329 92.5005
R1435 VDD.n5326 VDD.n5325 92.5005
R1436 VDD.n5322 VDD.n5321 92.5005
R1437 VDD.n5318 VDD.n5317 92.5005
R1438 VDD.n5314 VDD.n5313 92.5005
R1439 VDD.n5310 VDD.n5309 92.5005
R1440 VDD.n5306 VDD.n5305 92.5005
R1441 VDD.n5302 VDD.n5301 92.5005
R1442 VDD.n5298 VDD.n5297 92.5005
R1443 VDD.n5294 VDD.n5293 92.5005
R1444 VDD.n5290 VDD.n5289 92.5005
R1445 VDD.n5286 VDD.n5285 92.5005
R1446 VDD.n5282 VDD.n5281 92.5005
R1447 VDD.n13 VDD.n12 92.5005
R1448 VDD.n17 VDD.n16 92.5005
R1449 VDD.n21 VDD.n20 92.5005
R1450 VDD.n25 VDD.n24 92.5005
R1451 VDD.n29 VDD.n28 92.5005
R1452 VDD.n33 VDD.n32 92.5005
R1453 VDD.n37 VDD.n36 92.5005
R1454 VDD.n41 VDD.n40 92.5005
R1455 VDD.n45 VDD.n44 92.5005
R1456 VDD.n49 VDD.n48 92.5005
R1457 VDD.n53 VDD.n52 92.5005
R1458 VDD.n57 VDD.n56 92.5005
R1459 VDD.n61 VDD.n60 92.5005
R1460 VDD.n65 VDD.n64 92.5005
R1461 VDD.n69 VDD.n68 92.5005
R1462 VDD.n71 VDD.n70 92.5005
R1463 VDD.n73 VDD.n72 92.5005
R1464 VDD.n75 VDD.n74 92.5005
R1465 VDD.n6497 VDD.n6496 92.5005
R1466 VDD.n6495 VDD.n6494 92.5005
R1467 VDD.n5196 VDD.n5159 84.4449
R1468 VDD.n369 VDD.n368 69.3656
R1469 VDD.n5261 VDD.n5202 67.9542
R1470 VDD.n5261 VDD.n5203 67.9542
R1471 VDD.n5261 VDD.n5204 67.9542
R1472 VDD.n5261 VDD.n5205 67.9542
R1473 VDD.n5261 VDD.n5206 67.9542
R1474 VDD.n5261 VDD.n5207 67.9542
R1475 VDD.n5261 VDD.n5208 67.9542
R1476 VDD.n5261 VDD.n5209 67.9542
R1477 VDD.n5261 VDD.n5210 67.9542
R1478 VDD.n5261 VDD.n5211 67.9542
R1479 VDD.n5261 VDD.n5212 67.9542
R1480 VDD.n5261 VDD.n5213 67.9542
R1481 VDD.n5261 VDD.n5214 67.9542
R1482 VDD.n5261 VDD.n5215 67.9542
R1483 VDD.n5261 VDD.n5216 67.9542
R1484 VDD.n5261 VDD.n5217 67.9542
R1485 VDD.n5261 VDD.n5218 67.9542
R1486 VDD.n5261 VDD.n5219 67.9542
R1487 VDD.n5261 VDD.n5220 67.9542
R1488 VDD.n5261 VDD.n5221 67.9542
R1489 VDD.n5261 VDD.n5222 67.9542
R1490 VDD.n5261 VDD.n5223 67.9542
R1491 VDD.n5261 VDD.n5224 67.9542
R1492 VDD.n5261 VDD.n5225 67.9542
R1493 VDD.n5261 VDD.n5226 67.9542
R1494 VDD.n5261 VDD.n5227 67.9542
R1495 VDD.n5261 VDD.n5228 67.9542
R1496 VDD.n5261 VDD.n5229 67.9542
R1497 VDD.n5261 VDD.n5230 67.9542
R1498 VDD.n5261 VDD.n5235 67.9542
R1499 VDD.n5261 VDD.n5236 67.9542
R1500 VDD.n5261 VDD.n5237 67.9542
R1501 VDD.n5261 VDD.n5238 67.9542
R1502 VDD.n5261 VDD.n5239 67.9542
R1503 VDD.n5261 VDD.n5240 67.9542
R1504 VDD.n5261 VDD.n5241 67.9542
R1505 VDD.n5261 VDD.n5242 67.9542
R1506 VDD.n5261 VDD.n5243 67.9542
R1507 VDD.n5261 VDD.n5244 67.9542
R1508 VDD.n5261 VDD.n5245 67.9542
R1509 VDD.n5261 VDD.n5246 67.9542
R1510 VDD.n5261 VDD.n5247 67.9542
R1511 VDD.n5261 VDD.n5248 67.9542
R1512 VDD.n5261 VDD.n5249 67.9542
R1513 VDD.n5261 VDD.n5250 67.9542
R1514 VDD.n5261 VDD.n5251 67.9542
R1515 VDD.n5261 VDD.n5252 67.9542
R1516 VDD.n5261 VDD.n5253 67.9542
R1517 VDD.n5261 VDD.n5254 67.9542
R1518 VDD.n5261 VDD.n5255 67.9542
R1519 VDD.n5261 VDD.n5256 67.9542
R1520 VDD.n5261 VDD.n5257 67.9542
R1521 VDD.n5261 VDD.n5258 67.9542
R1522 VDD.n5261 VDD.n5259 67.9542
R1523 VDD.n1089 VDD.n1088 66.8854
R1524 VDD.n872 VDD.n871 66.3497
R1525 VDD.n1432 VDD.n1431 49.0945
R1526 VDD.n1435 VDD.n1434 49.0945
R1527 VDD.n1438 VDD.n1437 49.0945
R1528 VDD.n866 VDD.n865 44.768
R1529 VDD.n1305 VDD.t35 44.6138
R1530 VDD.n1443 VDD.n1442 41.6217
R1531 VDD.n5261 VDD.n5231 41.6217
R1532 VDD.n5261 VDD.n5260 41.6217
R1533 VDD.n1442 VDD.n1441 41.6215
R1534 VDD.n5261 VDD.n5201 41.6215
R1535 VDD.n5261 VDD.n5234 41.6215
R1536 VDD.n2986 VDD.n2985 38.7994
R1537 VDD.n1562 VDD.n1561 38.7994
R1538 VDD.n1544 VDD.n1543 38.7994
R1539 VDD.n1678 VDD.n1677 38.7994
R1540 VDD.n1700 VDD.n1699 38.7994
R1541 VDD.n1243 VDD.n1242 38.7994
R1542 VDD.n1427 VDD.n1426 38.7994
R1543 VDD.n1370 VDD.n1369 38.7994
R1544 VDD.n2986 VDD.n2984 38.7989
R1545 VDD.n1570 VDD.n1569 38.7989
R1546 VDD.n1552 VDD.n1551 38.7989
R1547 VDD.n1686 VDD.n1685 38.7989
R1548 VDD.n1708 VDD.n1707 38.7989
R1549 VDD.n1251 VDD.n1250 38.7989
R1550 VDD.n2983 VDD.n2981 38.7987
R1551 VDD.n2980 VDD.n2978 38.7987
R1552 VDD.n2977 VDD.n2975 38.7987
R1553 VDD.n2974 VDD.n2972 38.7987
R1554 VDD.n2971 VDD.n2969 38.7987
R1555 VDD.n2968 VDD.n2966 38.7987
R1556 VDD.n2965 VDD.n2963 38.7987
R1557 VDD.n2962 VDD.n2960 38.7987
R1558 VDD.n2959 VDD.n2957 38.7987
R1559 VDD.n2956 VDD.n2954 38.7987
R1560 VDD.n2953 VDD.n2951 38.7987
R1561 VDD.n2950 VDD.n2948 38.7987
R1562 VDD.n2947 VDD.n2945 38.7987
R1563 VDD.n2944 VDD.n2942 38.7987
R1564 VDD.n2983 VDD.n2982 38.7987
R1565 VDD.n2980 VDD.n2979 38.7987
R1566 VDD.n2977 VDD.n2976 38.7987
R1567 VDD.n2974 VDD.n2973 38.7987
R1568 VDD.n2971 VDD.n2970 38.7987
R1569 VDD.n2968 VDD.n2967 38.7987
R1570 VDD.n2965 VDD.n2964 38.7987
R1571 VDD.n2962 VDD.n2961 38.7987
R1572 VDD.n2959 VDD.n2958 38.7987
R1573 VDD.n2956 VDD.n2955 38.7987
R1574 VDD.n2953 VDD.n2952 38.7987
R1575 VDD.n2950 VDD.n2949 38.7987
R1576 VDD.n2947 VDD.n2946 38.7987
R1577 VDD.n2944 VDD.n2943 38.7987
R1578 VDD.n2941 VDD.n2940 38.7987
R1579 VDD.n2939 VDD.n2938 38.7987
R1580 VDD.n2937 VDD.n2935 38.7987
R1581 VDD.n2934 VDD.n2932 38.7987
R1582 VDD.n2931 VDD.n2929 38.7987
R1583 VDD.n2928 VDD.n2926 38.7987
R1584 VDD.n2925 VDD.n2923 38.7987
R1585 VDD.n2922 VDD.n2920 38.7987
R1586 VDD.n2919 VDD.n2917 38.7987
R1587 VDD.n2916 VDD.n2914 38.7987
R1588 VDD.n2913 VDD.n2911 38.7987
R1589 VDD.n2910 VDD.n2908 38.7987
R1590 VDD.n2907 VDD.n2905 38.7987
R1591 VDD.n2904 VDD.n2902 38.7987
R1592 VDD.n2937 VDD.n2936 38.7987
R1593 VDD.n2934 VDD.n2933 38.7987
R1594 VDD.n2931 VDD.n2930 38.7987
R1595 VDD.n2928 VDD.n2927 38.7987
R1596 VDD.n2925 VDD.n2924 38.7987
R1597 VDD.n2922 VDD.n2921 38.7987
R1598 VDD.n2919 VDD.n2918 38.7987
R1599 VDD.n2916 VDD.n2915 38.7987
R1600 VDD.n2913 VDD.n2912 38.7987
R1601 VDD.n2910 VDD.n2909 38.7987
R1602 VDD.n2907 VDD.n2906 38.7987
R1603 VDD.n2904 VDD.n2903 38.7987
R1604 VDD.n1233 VDD.n1232 38.7987
R1605 VDD.n1225 VDD.n1224 38.7987
R1606 VDD.n1421 VDD.n1420 38.7987
R1607 VDD.n1416 VDD.n1415 38.7987
R1608 VDD.n1364 VDD.n1363 38.7987
R1609 VDD.n1359 VDD.n1358 38.7987
R1610 VDD.n374 VDD.n373 34.4176
R1611 VDD.n875 VDD.n874 34.2738
R1612 VDD.n1085 VDD.n1082 33.4435
R1613 VDD.n1094 VDD.n1091 33.4435
R1614 VDD.n1089 VDD.n1087 33.4435
R1615 VDD.n1100 VDD.n1097 33.4435
R1616 VDD.n874 VDD.n870 33.4435
R1617 VDD.n373 VDD.n370 33.4435
R1618 VDD.n6488 VDD.n6486 33.4435
R1619 VDD.n6491 VDD.n6489 33.4435
R1620 VDD.n1100 VDD.n1099 33.4431
R1621 VDD.n1085 VDD.n1084 33.4431
R1622 VDD.n1094 VDD.n1093 33.4431
R1623 VDD.n874 VDD.n873 33.4431
R1624 VDD.n358 VDD.n357 33.4431
R1625 VDD.n373 VDD.n372 33.4431
R1626 VDD.n6488 VDD.n6487 33.4431
R1627 VDD.n6491 VDD.n6490 33.4431
R1628 VDD.n2839 VDD.n2838 33.4428
R1629 VDD.n2890 VDD.n2888 33.4428
R1630 VDD.n2887 VDD.n2885 33.4428
R1631 VDD.n2884 VDD.n2882 33.4428
R1632 VDD.n2881 VDD.n2879 33.4428
R1633 VDD.n2878 VDD.n2876 33.4428
R1634 VDD.n2875 VDD.n2873 33.4428
R1635 VDD.n2872 VDD.n2870 33.4428
R1636 VDD.n2890 VDD.n2889 33.4428
R1637 VDD.n2887 VDD.n2886 33.4428
R1638 VDD.n2884 VDD.n2883 33.4428
R1639 VDD.n2881 VDD.n2880 33.4428
R1640 VDD.n2878 VDD.n2877 33.4428
R1641 VDD.n2875 VDD.n2874 33.4428
R1642 VDD.n2872 VDD.n2871 33.4428
R1643 VDD.n2869 VDD.n2868 33.4428
R1644 VDD.n2841 VDD.n2840 33.4428
R1645 VDD.n2837 VDD.n2836 31.4488
R1646 VDD.n3029 VDD.n3028 31.4488
R1647 VDD.n3695 VDD.n3694 31.4488
R1648 VDD.n3716 VDD.n3715 31.4488
R1649 VDD.n4055 VDD.n4054 31.4488
R1650 VDD.n4072 VDD.n4071 31.4488
R1651 VDD.n4376 VDD.n4375 31.4488
R1652 VDD.n4393 VDD.n4392 31.4488
R1653 VDD.n4722 VDD.n4721 31.4488
R1654 VDD.n4741 VDD.n4740 31.4488
R1655 VDD.n5077 VDD.n5076 31.4488
R1656 VDD.n5092 VDD.n5091 31.4488
R1657 VDD.n1278 VDD.t37 30.1801
R1658 VDD.n1263 VDD.t39 30.1801
R1659 VDD.n1717 VDD.t446 30.1801
R1660 VDD.n1734 VDD.t452 30.1801
R1661 VDD.n1759 VDD.t31 30.1801
R1662 VDD.n1777 VDD.t140 30.1801
R1663 VDD.n1651 VDD.t159 30.1801
R1664 VDD.n1633 VDD.t161 30.1801
R1665 VDD.n1608 VDD.t155 30.1801
R1666 VDD.n1590 VDD.t157 30.1801
R1667 VDD.n1448 VDD.t59 30.1801
R1668 VDD.n1463 VDD.t57 30.1801
R1669 VDD.n1483 VDD.t53 30.1801
R1670 VDD.n1498 VDD.t55 30.1801
R1671 VDD.n1255 VDD.n1252 30.1181
R1672 VDD.n1747 VDD.n1709 30.1181
R1673 VDD.n1694 VDD.n1691 30.1181
R1674 VDD.n1790 VDD.n1687 30.1181
R1675 VDD.n1672 VDD.n1669 30.1181
R1676 VDD.n1621 VDD.n1553 30.1181
R1677 VDD.n1538 VDD.n1535 30.1181
R1678 VDD.n1579 VDD.n1571 30.1181
R1679 VDD.n1290 VDD.n1234 30.1181
R1680 VDD.n1347 VDD.n1325 30.1181
R1681 VDD.n1473 VDD.n1445 30.1181
R1682 VDD.n1400 VDD.n1381 30.1181
R1683 VDD.n1444 VDD.n1443 30.0704
R1684 VDD.n2693 VDD.n2692 29.5303
R1685 VDD.n1103 VDD.n1094 29.5303
R1686 VDD.n1103 VDD.n1089 29.5303
R1687 VDD.n1103 VDD.n1100 29.5303
R1688 VDD.n1103 VDD.n1085 29.5303
R1689 VDD.n357 VDD.n356 29.5303
R1690 VDD.n5195 VDD.n5194 29.5303
R1691 VDD.n5195 VDD.n5193 29.5303
R1692 VDD.n5195 VDD.n5192 29.5303
R1693 VDD.n5195 VDD.n5191 29.5303
R1694 VDD.n5195 VDD.n5190 29.5303
R1695 VDD.n5195 VDD.n5189 29.5303
R1696 VDD.n5195 VDD.n5188 29.5303
R1697 VDD.n5195 VDD.n5187 29.5303
R1698 VDD.n5195 VDD.n5186 29.5303
R1699 VDD.n5195 VDD.n5185 29.5303
R1700 VDD.n5195 VDD.n5184 29.5303
R1701 VDD.n5195 VDD.n5183 29.5303
R1702 VDD.n5195 VDD.n5182 29.5303
R1703 VDD.n5195 VDD.n5181 29.5303
R1704 VDD.n5195 VDD.n5180 29.5303
R1705 VDD.n5195 VDD.n5179 29.5303
R1706 VDD.n5195 VDD.n5178 29.5303
R1707 VDD.n5195 VDD.n5177 29.5303
R1708 VDD.n5195 VDD.n5176 29.5303
R1709 VDD.n5195 VDD.n5175 29.5303
R1710 VDD.n5195 VDD.n5174 29.5303
R1711 VDD.n5195 VDD.n5173 29.5303
R1712 VDD.n5195 VDD.n5172 29.5303
R1713 VDD.n5195 VDD.n5171 29.5303
R1714 VDD.n5195 VDD.n5170 29.5303
R1715 VDD.n5195 VDD.n5169 29.5303
R1716 VDD.n5195 VDD.n5168 29.5303
R1717 VDD.n5195 VDD.n5167 29.5303
R1718 VDD.n5195 VDD.n5166 29.5303
R1719 VDD.n5195 VDD.n5165 29.5303
R1720 VDD.n5195 VDD.n5164 29.5303
R1721 VDD.n5195 VDD.n5163 29.5303
R1722 VDD.n5195 VDD.n5162 29.5303
R1723 VDD.n5195 VDD.n5161 29.5303
R1724 VDD.n5195 VDD.n5160 29.5303
R1725 VDD.n6492 VDD.n6488 29.5303
R1726 VDD.n6492 VDD.n6491 29.5303
R1727 VDD.n2891 VDD.n2890 29.5301
R1728 VDD.n2891 VDD.n2887 29.5301
R1729 VDD.n2891 VDD.n2884 29.5301
R1730 VDD.n2891 VDD.n2881 29.5301
R1731 VDD.n2891 VDD.n2878 29.5301
R1732 VDD.n2891 VDD.n2875 29.5301
R1733 VDD.n2891 VDD.n2872 29.5301
R1734 VDD.n2891 VDD.n2869 29.5301
R1735 VDD.n2891 VDD.n2867 29.5301
R1736 VDD.n2891 VDD.n2866 29.5301
R1737 VDD.n2891 VDD.n2865 29.5301
R1738 VDD.n2891 VDD.n2864 29.5301
R1739 VDD.n2891 VDD.n2863 29.5301
R1740 VDD.n2891 VDD.n2862 29.5301
R1741 VDD.n2891 VDD.n2861 29.5301
R1742 VDD.n2891 VDD.n2860 29.5301
R1743 VDD.n2891 VDD.n2859 29.5301
R1744 VDD.n2891 VDD.n2858 29.5301
R1745 VDD.n2891 VDD.n2857 29.5301
R1746 VDD.n2891 VDD.n2856 29.5301
R1747 VDD.n2891 VDD.n2855 29.5301
R1748 VDD.n2891 VDD.n2854 29.5301
R1749 VDD.n2891 VDD.n2853 29.5301
R1750 VDD.n2891 VDD.n2852 29.5301
R1751 VDD.n2891 VDD.n2851 29.5301
R1752 VDD.n2891 VDD.n2850 29.5301
R1753 VDD.n2891 VDD.n2849 29.5301
R1754 VDD.n2891 VDD.n2848 29.5301
R1755 VDD.n2891 VDD.n2847 29.5301
R1756 VDD.n2891 VDD.n2846 29.5301
R1757 VDD.n2891 VDD.n2845 29.5301
R1758 VDD.n2891 VDD.n2844 29.5301
R1759 VDD.n2891 VDD.n2843 29.5301
R1760 VDD.n2891 VDD.n2842 29.5301
R1761 VDD.n2891 VDD.n2841 29.5301
R1762 VDD.n2891 VDD.n2839 29.5301
R1763 VDD.n3509 VDD.n3498 29.4833
R1764 VDD.n3553 VDD.n3542 29.4833
R1765 VDD.n3875 VDD.n3862 29.4833
R1766 VDD.n3914 VDD.n3905 29.4833
R1767 VDD.n4213 VDD.n4207 29.4833
R1768 VDD.n4248 VDD.n4241 29.4833
R1769 VDD.n4543 VDD.n4534 29.4833
R1770 VDD.n4580 VDD.n4569 29.4833
R1771 VDD.n4897 VDD.n4886 29.4833
R1772 VDD.n4936 VDD.n4925 29.4833
R1773 VDD.n6210 VDD.t7 27.6955
R1774 VDD.n6210 VDD.t450 27.6955
R1775 VDD.n6203 VDD.t43 27.6955
R1776 VDD.n6203 VDD.t101 27.6955
R1777 VDD.n6196 VDD.t460 27.6955
R1778 VDD.n6196 VDD.t462 27.6955
R1779 VDD.n6189 VDD.t383 27.6955
R1780 VDD.n6189 VDD.t151 27.6955
R1781 VDD.n6182 VDD.t398 27.6955
R1782 VDD.n6182 VDD.t82 27.6955
R1783 VDD.n6175 VDD.t10 27.6955
R1784 VDD.n6175 VDD.t20 27.6955
R1785 VDD.n6168 VDD.t137 27.6955
R1786 VDD.n6168 VDD.t87 27.6955
R1787 VDD.n6161 VDD.t73 27.6955
R1788 VDD.n6161 VDD.t48 27.6955
R1789 VDD.n6154 VDD.t136 27.6955
R1790 VDD.n6154 VDD.t376 27.6955
R1791 VDD.n6147 VDD.t464 27.6955
R1792 VDD.n6147 VDD.t463 27.6955
R1793 VDD.n6140 VDD.t393 27.6955
R1794 VDD.n6140 VDD.t131 27.6955
R1795 VDD.n6133 VDD.t122 27.6955
R1796 VDD.n6133 VDD.t384 27.6955
R1797 VDD.n6126 VDD.t97 27.6955
R1798 VDD.n6126 VDD.t371 27.6955
R1799 VDD.n6119 VDD.t372 27.6955
R1800 VDD.n6119 VDD.t107 27.6955
R1801 VDD.n6112 VDD.t387 27.6955
R1802 VDD.n6112 VDD.t449 27.6955
R1803 VDD.n6105 VDD.t16 27.6955
R1804 VDD.n6105 VDD.t9 27.6955
R1805 VDD.n6098 VDD.t3 27.6955
R1806 VDD.n6098 VDD.t413 27.6955
R1807 VDD.n6091 VDD.t104 27.6955
R1808 VDD.n6091 VDD.t139 27.6955
R1809 VDD.n6084 VDD.t459 27.6955
R1810 VDD.n6084 VDD.t381 27.6955
R1811 VDD.n6077 VDD.t121 27.6955
R1812 VDD.n6077 VDD.t385 27.6955
R1813 VDD.n6031 VDD.t424 27.6955
R1814 VDD.n6031 VDD.t62 27.6955
R1815 VDD.n6024 VDD.t400 27.6955
R1816 VDD.n6024 VDD.t103 27.6955
R1817 VDD.n6017 VDD.t89 27.6955
R1818 VDD.n6017 VDD.t396 27.6955
R1819 VDD.n6010 VDD.t369 27.6955
R1820 VDD.n6010 VDD.t149 27.6955
R1821 VDD.n6003 VDD.t124 27.6955
R1822 VDD.n6003 VDD.t432 27.6955
R1823 VDD.n5996 VDD.t1 27.6955
R1824 VDD.n5996 VDD.t453 27.6955
R1825 VDD.n5989 VDD.t166 27.6955
R1826 VDD.n5989 VDD.t410 27.6955
R1827 VDD.n5982 VDD.t439 27.6955
R1828 VDD.n5982 VDD.t433 27.6955
R1829 VDD.n5975 VDD.t150 27.6955
R1830 VDD.n5975 VDD.t134 27.6955
R1831 VDD.n5968 VDD.t69 27.6955
R1832 VDD.n5968 VDD.t106 27.6955
R1833 VDD.n5961 VDD.t145 27.6955
R1834 VDD.n5961 VDD.t154 27.6955
R1835 VDD.n5954 VDD.t85 27.6955
R1836 VDD.n5954 VDD.t90 27.6955
R1837 VDD.n5947 VDD.t390 27.6955
R1838 VDD.n5947 VDD.t111 27.6955
R1839 VDD.n5940 VDD.t51 27.6955
R1840 VDD.n5940 VDD.t427 27.6955
R1841 VDD.n5933 VDD.t377 27.6955
R1842 VDD.n5933 VDD.t94 27.6955
R1843 VDD.n5926 VDD.t379 27.6955
R1844 VDD.n5926 VDD.t426 27.6955
R1845 VDD.n5919 VDD.t454 27.6955
R1846 VDD.n5919 VDD.t420 27.6955
R1847 VDD.n5912 VDD.t438 27.6955
R1848 VDD.n5912 VDD.t457 27.6955
R1849 VDD.n5905 VDD.t392 27.6955
R1850 VDD.n5905 VDD.t125 27.6955
R1851 VDD.n5898 VDD.t447 27.6955
R1852 VDD.n5898 VDD.t32 27.6955
R1853 VDD.n5852 VDD.t402 27.6955
R1854 VDD.n5852 VDD.t448 27.6955
R1855 VDD.n5845 VDD.t403 27.6955
R1856 VDD.n5845 VDD.t46 27.6955
R1857 VDD.n5838 VDD.t132 27.6955
R1858 VDD.n5838 VDD.t30 27.6955
R1859 VDD.n5831 VDD.t373 27.6955
R1860 VDD.n5831 VDD.t407 27.6955
R1861 VDD.n5824 VDD.t401 27.6955
R1862 VDD.n5824 VDD.t64 27.6955
R1863 VDD.n5817 VDD.t67 27.6955
R1864 VDD.n5817 VDD.t429 27.6955
R1865 VDD.n5810 VDD.t113 27.6955
R1866 VDD.n5810 VDD.t126 27.6955
R1867 VDD.n5803 VDD.t374 27.6955
R1868 VDD.n5803 VDD.t65 27.6955
R1869 VDD.n5796 VDD.t445 27.6955
R1870 VDD.n5796 VDD.t421 27.6955
R1871 VDD.n5789 VDD.t119 27.6955
R1872 VDD.n5789 VDD.t147 27.6955
R1873 VDD.n5782 VDD.t416 27.6955
R1874 VDD.n5782 VDD.t130 27.6955
R1875 VDD.n5775 VDD.t102 27.6955
R1876 VDD.n5775 VDD.t409 27.6955
R1877 VDD.n5768 VDD.t434 27.6955
R1878 VDD.n5768 VDD.t123 27.6955
R1879 VDD.n5761 VDD.t66 27.6955
R1880 VDD.n5761 VDD.t148 27.6955
R1881 VDD.n5754 VDD.t116 27.6955
R1882 VDD.n5754 VDD.t114 27.6955
R1883 VDD.n5747 VDD.t437 27.6955
R1884 VDD.n5747 VDD.t112 27.6955
R1885 VDD.n5740 VDD.t406 27.6955
R1886 VDD.n5740 VDD.t388 27.6955
R1887 VDD.n5733 VDD.t164 27.6955
R1888 VDD.n5733 VDD.t382 27.6955
R1889 VDD.n5726 VDD.t418 27.6955
R1890 VDD.n5726 VDD.t118 27.6955
R1891 VDD.n5719 VDD.t441 27.6955
R1892 VDD.n5719 VDD.t108 27.6955
R1893 VDD.n5673 VDD.t430 27.6955
R1894 VDD.n5673 VDD.t440 27.6955
R1895 VDD.n5666 VDD.t44 27.6955
R1896 VDD.n5666 VDD.t146 27.6955
R1897 VDD.n5659 VDD.t386 27.6955
R1898 VDD.n5659 VDD.t442 27.6955
R1899 VDD.n5652 VDD.t425 27.6955
R1900 VDD.n5652 VDD.t144 27.6955
R1901 VDD.n5645 VDD.t86 27.6955
R1902 VDD.n5645 VDD.t5 27.6955
R1903 VDD.n5638 VDD.t41 27.6955
R1904 VDD.n5638 VDD.t138 27.6955
R1905 VDD.n5631 VDD.t92 27.6955
R1906 VDD.n5631 VDD.t12 27.6955
R1907 VDD.n5624 VDD.t404 27.6955
R1908 VDD.n5624 VDD.t49 27.6955
R1909 VDD.n5617 VDD.t451 27.6955
R1910 VDD.n5617 VDD.t370 27.6955
R1911 VDD.n5610 VDD.t34 27.6955
R1912 VDD.n5610 VDD.t375 27.6955
R1913 VDD.n5603 VDD.t26 27.6955
R1914 VDD.n5603 VDD.t417 27.6955
R1915 VDD.n5596 VDD.t455 27.6955
R1916 VDD.n5596 VDD.t28 27.6955
R1917 VDD.n5589 VDD.t75 27.6955
R1918 VDD.n5589 VDD.t431 27.6955
R1919 VDD.n5582 VDD.t395 27.6955
R1920 VDD.n5582 VDD.t95 27.6955
R1921 VDD.n5575 VDD.t399 27.6955
R1922 VDD.n5575 VDD.t96 27.6955
R1923 VDD.n5568 VDD.t109 27.6955
R1924 VDD.n5568 VDD.t415 27.6955
R1925 VDD.n5561 VDD.t74 27.6955
R1926 VDD.n5561 VDD.t412 27.6955
R1927 VDD.n5554 VDD.t84 27.6955
R1928 VDD.n5554 VDD.t163 27.6955
R1929 VDD.n5547 VDD.t77 27.6955
R1930 VDD.n5547 VDD.t422 27.6955
R1931 VDD.n5540 VDD.t128 27.6955
R1932 VDD.n5540 VDD.t25 27.6955
R1933 VDD.n5494 VDD.t456 27.6955
R1934 VDD.n5494 VDD.t414 27.6955
R1935 VDD.n5487 VDD.t165 27.6955
R1936 VDD.n5487 VDD.t458 27.6955
R1937 VDD.n5480 VDD.t436 27.6955
R1938 VDD.n5480 VDD.t100 27.6955
R1939 VDD.n5473 VDD.t18 27.6955
R1940 VDD.n5473 VDD.t397 27.6955
R1941 VDD.n5466 VDD.t81 27.6955
R1942 VDD.n5466 VDD.t391 27.6955
R1943 VDD.n5459 VDD.t435 27.6955
R1944 VDD.n5459 VDD.t152 27.6955
R1945 VDD.n5452 VDD.t444 27.6955
R1946 VDD.n5452 VDD.t127 27.6955
R1947 VDD.n5445 VDD.t419 27.6955
R1948 VDD.n5445 VDD.t141 27.6955
R1949 VDD.n5438 VDD.t461 27.6955
R1950 VDD.n5438 VDD.t423 27.6955
R1951 VDD.n5431 VDD.t142 27.6955
R1952 VDD.n5431 VDD.t167 27.6955
R1953 VDD.n5424 VDD.t14 27.6955
R1954 VDD.n5424 VDD.t466 27.6955
R1955 VDD.n5417 VDD.t79 27.6955
R1956 VDD.n5417 VDD.t153 27.6955
R1957 VDD.n5410 VDD.t71 27.6955
R1958 VDD.n5410 VDD.t428 27.6955
R1959 VDD.n5403 VDD.t465 27.6955
R1960 VDD.n5403 VDD.t22 27.6955
R1961 VDD.n5396 VDD.t394 27.6955
R1962 VDD.n5396 VDD.t405 27.6955
R1963 VDD.n5389 VDD.t52 27.6955
R1964 VDD.n5389 VDD.t68 27.6955
R1965 VDD.n5382 VDD.t378 27.6955
R1966 VDD.n5382 VDD.t408 27.6955
R1967 VDD.n5375 VDD.t443 27.6955
R1968 VDD.n5375 VDD.t99 27.6955
R1969 VDD.n5368 VDD.t411 27.6955
R1970 VDD.n5368 VDD.t389 27.6955
R1971 VDD.n5361 VDD.t380 27.6955
R1972 VDD.n5361 VDD.t63 27.6955
R1973 VDD.n2646 VDD.t229 27.6955
R1974 VDD.n2646 VDD.t327 27.6955
R1975 VDD.n2639 VDD.t238 27.6955
R1976 VDD.n2639 VDD.t337 27.6955
R1977 VDD.n2632 VDD.t326 27.6955
R1978 VDD.n2632 VDD.t175 27.6955
R1979 VDD.n2625 VDD.t258 27.6955
R1980 VDD.n2625 VDD.t306 27.6955
R1981 VDD.n2618 VDD.t207 27.6955
R1982 VDD.n2618 VDD.t197 27.6955
R1983 VDD.n2611 VDD.t280 27.6955
R1984 VDD.n2611 VDD.t335 27.6955
R1985 VDD.n2604 VDD.t184 27.6955
R1986 VDD.n2604 VDD.t263 27.6955
R1987 VDD.n2597 VDD.t329 27.6955
R1988 VDD.n2597 VDD.t202 27.6955
R1989 VDD.n2590 VDD.t358 27.6955
R1990 VDD.n2590 VDD.t308 27.6955
R1991 VDD.n2583 VDD.t218 27.6955
R1992 VDD.n2583 VDD.t216 27.6955
R1993 VDD.n2576 VDD.t325 27.6955
R1994 VDD.n2576 VDD.t262 27.6955
R1995 VDD.n2569 VDD.t182 27.6955
R1996 VDD.n2569 VDD.t334 27.6955
R1997 VDD.n2562 VDD.t340 27.6955
R1998 VDD.n2562 VDD.t240 27.6955
R1999 VDD.n2555 VDD.t204 27.6955
R2000 VDD.n2555 VDD.t235 27.6955
R2001 VDD.n2548 VDD.t191 27.6955
R2002 VDD.n2548 VDD.t354 27.6955
R2003 VDD.n2541 VDD.t304 27.6955
R2004 VDD.n2541 VDD.t255 27.6955
R2005 VDD.n2534 VDD.t169 27.6955
R2006 VDD.n2534 VDD.t245 27.6955
R2007 VDD.n2527 VDD.t214 27.6955
R2008 VDD.n2527 VDD.t170 27.6955
R2009 VDD.n2520 VDD.t320 27.6955
R2010 VDD.n2520 VDD.t226 27.6955
R2011 VDD.n2513 VDD.t186 27.6955
R2012 VDD.n2513 VDD.t343 27.6955
R2013 VDD.n2467 VDD.t365 27.6955
R2014 VDD.n2467 VDD.t249 27.6955
R2015 VDD.n2460 VDD.t173 27.6955
R2016 VDD.n2460 VDD.t257 27.6955
R2017 VDD.n2453 VDD.t248 27.6955
R2018 VDD.n2453 VDD.t294 27.6955
R2019 VDD.n2446 VDD.t199 27.6955
R2020 VDD.n2446 VDD.t237 27.6955
R2021 VDD.n2439 VDD.t331 27.6955
R2022 VDD.n2439 VDD.t319 27.6955
R2023 VDD.n2432 VDD.t221 27.6955
R2024 VDD.n2432 VDD.t250 27.6955
R2025 VDD.n2425 VDD.t303 27.6955
R2026 VDD.n2425 VDD.t205 27.6955
R2027 VDD.n2418 VDD.t251 27.6955
R2028 VDD.n2418 VDD.t324 27.6955
R2029 VDD.n2411 VDD.t275 27.6955
R2030 VDD.n2411 VDD.t236 27.6955
R2031 VDD.n2404 VDD.t344 27.6955
R2032 VDD.n2404 VDD.t355 27.6955
R2033 VDD.n2397 VDD.t247 27.6955
R2034 VDD.n2397 VDD.t203 27.6955
R2035 VDD.n2390 VDD.t302 27.6955
R2036 VDD.n2390 VDD.t254 27.6955
R2037 VDD.n2383 VDD.t259 27.6955
R2038 VDD.n2383 VDD.t177 27.6955
R2039 VDD.n2376 VDD.t330 27.6955
R2040 VDD.n2376 VDD.t168 27.6955
R2041 VDD.n2369 VDD.t318 27.6955
R2042 VDD.n2369 VDD.t271 27.6955
R2043 VDD.n2362 VDD.t232 27.6955
R2044 VDD.n2362 VDD.t195 27.6955
R2045 VDD.n2355 VDD.t288 27.6955
R2046 VDD.n2355 VDD.t188 27.6955
R2047 VDD.n2348 VDD.t342 27.6955
R2048 VDD.n2348 VDD.t290 27.6955
R2049 VDD.n2341 VDD.t244 27.6955
R2050 VDD.n2341 VDD.t361 27.6955
R2051 VDD.n2334 VDD.t310 27.6955
R2052 VDD.n2334 VDD.t261 27.6955
R2053 VDD.n2288 VDD.t212 27.6955
R2054 VDD.n2288 VDD.t299 27.6955
R2055 VDD.n2281 VDD.t219 27.6955
R2056 VDD.n2281 VDD.t309 27.6955
R2057 VDD.n2274 VDD.t296 27.6955
R2058 VDD.n2274 VDD.t350 27.6955
R2059 VDD.n2267 VDD.t239 27.6955
R2060 VDD.n2267 VDD.t279 27.6955
R2061 VDD.n2260 VDD.t180 27.6955
R2062 VDD.n2260 VDD.t172 27.6955
R2063 VDD.n2253 VDD.t256 27.6955
R2064 VDD.n2253 VDD.t307 27.6955
R2065 VDD.n2246 VDD.t357 27.6955
R2066 VDD.n2246 VDD.t242 27.6955
R2067 VDD.n2239 VDD.t300 27.6955
R2068 VDD.n2239 VDD.t176 27.6955
R2069 VDD.n2232 VDD.t328 27.6955
R2070 VDD.n2232 VDD.t276 27.6955
R2071 VDD.n2225 VDD.t193 27.6955
R2072 VDD.n2225 VDD.t201 27.6955
R2073 VDD.n2218 VDD.t295 27.6955
R2074 VDD.n2218 VDD.t241 27.6955
R2075 VDD.n2211 VDD.t356 27.6955
R2076 VDD.n2211 VDD.t305 27.6955
R2077 VDD.n2204 VDD.t312 27.6955
R2078 VDD.n2204 VDD.t222 27.6955
R2079 VDD.n2197 VDD.t179 27.6955
R2080 VDD.n2197 VDD.t217 27.6955
R2081 VDD.n2190 VDD.t171 27.6955
R2082 VDD.n2190 VDD.t321 27.6955
R2083 VDD.n2183 VDD.t272 27.6955
R2084 VDD.n2183 VDD.t233 27.6955
R2085 VDD.n2176 VDD.t345 27.6955
R2086 VDD.n2176 VDD.t227 27.6955
R2087 VDD.n2169 VDD.t190 27.6955
R2088 VDD.n2169 VDD.t346 27.6955
R2089 VDD.n2162 VDD.t291 27.6955
R2090 VDD.n2162 VDD.t208 27.6955
R2091 VDD.n2155 VDD.t362 27.6955
R2092 VDD.n2155 VDD.t313 27.6955
R2093 VDD.n2112 VDD.t200 27.6955
R2094 VDD.n2112 VDD.t285 27.6955
R2095 VDD.n2105 VDD.t209 27.6955
R2096 VDD.n2105 VDD.t292 27.6955
R2097 VDD.n2098 VDD.t284 27.6955
R2098 VDD.n2098 VDD.t338 27.6955
R2099 VDD.n2091 VDD.t228 27.6955
R2100 VDD.n2091 VDD.t266 27.6955
R2101 VDD.n2084 VDD.t367 27.6955
R2102 VDD.n2084 VDD.t360 27.6955
R2103 VDD.n2077 VDD.t243 27.6955
R2104 VDD.n2077 VDD.t289 27.6955
R2105 VDD.n2070 VDD.t341 27.6955
R2106 VDD.n2070 VDD.t231 27.6955
R2107 VDD.n2063 VDD.t286 27.6955
R2108 VDD.n2063 VDD.t363 27.6955
R2109 VDD.n2056 VDD.t315 27.6955
R2110 VDD.n2056 VDD.t264 27.6955
R2111 VDD.n2049 VDD.t181 27.6955
R2112 VDD.n2049 VDD.t189 27.6955
R2113 VDD.n2042 VDD.t282 27.6955
R2114 VDD.n2042 VDD.t230 27.6955
R2115 VDD.n2035 VDD.t339 27.6955
R2116 VDD.n2035 VDD.t287 27.6955
R2117 VDD.n2028 VDD.t298 27.6955
R2118 VDD.n2028 VDD.t211 27.6955
R2119 VDD.n2021 VDD.t366 27.6955
R2120 VDD.n2021 VDD.t206 27.6955
R2121 VDD.n2014 VDD.t359 27.6955
R2122 VDD.n2014 VDD.t311 27.6955
R2123 VDD.n2007 VDD.t260 27.6955
R2124 VDD.n2007 VDD.t225 27.6955
R2125 VDD.n2000 VDD.t332 27.6955
R2126 VDD.n2000 VDD.t215 27.6955
R2127 VDD.n1993 VDD.t178 27.6955
R2128 VDD.n1993 VDD.t333 27.6955
R2129 VDD.n1986 VDD.t278 27.6955
R2130 VDD.n1986 VDD.t196 27.6955
R2131 VDD.n1979 VDD.t349 27.6955
R2132 VDD.n1979 VDD.t301 27.6955
R2133 VDD.n1933 VDD.t185 27.6955
R2134 VDD.n1933 VDD.t269 27.6955
R2135 VDD.n1926 VDD.t194 27.6955
R2136 VDD.n1926 VDD.t277 27.6955
R2137 VDD.n1919 VDD.t268 27.6955
R2138 VDD.n1919 VDD.t317 27.6955
R2139 VDD.n1912 VDD.t220 27.6955
R2140 VDD.n1912 VDD.t253 27.6955
R2141 VDD.n1905 VDD.t353 27.6955
R2142 VDD.n1905 VDD.t348 27.6955
R2143 VDD.n1898 VDD.t234 27.6955
R2144 VDD.n1898 VDD.t274 27.6955
R2145 VDD.n1891 VDD.t323 27.6955
R2146 VDD.n1891 VDD.t224 27.6955
R2147 VDD.n1884 VDD.t270 27.6955
R2148 VDD.n1884 VDD.t351 27.6955
R2149 VDD.n1877 VDD.t297 27.6955
R2150 VDD.n1877 VDD.t252 27.6955
R2151 VDD.n1870 VDD.t368 27.6955
R2152 VDD.n1870 VDD.t174 27.6955
R2153 VDD.n1863 VDD.t267 27.6955
R2154 VDD.n1863 VDD.t223 27.6955
R2155 VDD.n1856 VDD.t322 27.6955
R2156 VDD.n1856 VDD.t273 27.6955
R2157 VDD.n1849 VDD.t281 27.6955
R2158 VDD.n1849 VDD.t198 27.6955
R2159 VDD.n1842 VDD.t352 27.6955
R2160 VDD.n1842 VDD.t192 27.6955
R2161 VDD.n1835 VDD.t347 27.6955
R2162 VDD.n1835 VDD.t293 27.6955
R2163 VDD.n1828 VDD.t246 27.6955
R2164 VDD.n1828 VDD.t213 27.6955
R2165 VDD.n1821 VDD.t314 27.6955
R2166 VDD.n1821 VDD.t210 27.6955
R2167 VDD.n1814 VDD.t364 27.6955
R2168 VDD.n1814 VDD.t316 27.6955
R2169 VDD.n1807 VDD.t265 27.6955
R2170 VDD.n1807 VDD.t183 27.6955
R2171 VDD.n1800 VDD.t336 27.6955
R2172 VDD.n1800 VDD.t283 27.6955
R2173 VDD.n106 VDD.t36 27.6955
R2174 VDD.n1378 VDD.t54 27.6955
R2175 VDD.n1378 VDD.t56 27.6955
R2176 VDD.n1377 VDD.t60 27.6955
R2177 VDD.n1377 VDD.t58 27.6955
R2178 VDD.n1376 VDD.t156 27.6955
R2179 VDD.n1376 VDD.t158 27.6955
R2180 VDD.n1375 VDD.t160 27.6955
R2181 VDD.n1375 VDD.t162 27.6955
R2182 VDD.n1209 VDD.t38 27.6955
R2183 VDD.n1209 VDD.t40 27.6955
R2184 VDD.n3008 VDD.n3007 27.5177
R2185 VDD.n3672 VDD.n3671 27.5177
R2186 VDD.n3735 VDD.n3734 27.5177
R2187 VDD.n4035 VDD.n4034 27.5177
R2188 VDD.n4090 VDD.n4089 27.5177
R2189 VDD.n4358 VDD.n4357 27.5177
R2190 VDD.n4412 VDD.n4411 27.5177
R2191 VDD.n4702 VDD.n4701 27.5177
R2192 VDD.n4760 VDD.n4759 27.5177
R2193 VDD.n5056 VDD.n5055 27.5177
R2194 VDD.n5111 VDD.n5110 27.5177
R2195 VDD.n2987 VDD.n2986 26.8524
R2196 VDD.n1568 VDD.n1567 26.8524
R2197 VDD.n1569 VDD.n1568 26.8524
R2198 VDD.n1550 VDD.n1549 26.8524
R2199 VDD.n1551 VDD.n1550 26.8524
R2200 VDD.n1684 VDD.n1683 26.8524
R2201 VDD.n1685 VDD.n1684 26.8524
R2202 VDD.n1706 VDD.n1705 26.8524
R2203 VDD.n1707 VDD.n1706 26.8524
R2204 VDD.n1249 VDD.n1248 26.8524
R2205 VDD.n1250 VDD.n1249 26.8524
R2206 VDD.n1426 VDD.n1425 26.8524
R2207 VDD.n1369 VDD.n1368 26.8524
R2208 VDD.n2987 VDD.n2983 26.8521
R2209 VDD.n2987 VDD.n2980 26.8521
R2210 VDD.n2987 VDD.n2977 26.8521
R2211 VDD.n2987 VDD.n2974 26.8521
R2212 VDD.n2987 VDD.n2971 26.8521
R2213 VDD.n2987 VDD.n2968 26.8521
R2214 VDD.n2987 VDD.n2965 26.8521
R2215 VDD.n2987 VDD.n2962 26.8521
R2216 VDD.n2987 VDD.n2959 26.8521
R2217 VDD.n2987 VDD.n2956 26.8521
R2218 VDD.n2987 VDD.n2953 26.8521
R2219 VDD.n2987 VDD.n2950 26.8521
R2220 VDD.n2987 VDD.n2947 26.8521
R2221 VDD.n2987 VDD.n2944 26.8521
R2222 VDD.n2987 VDD.n2941 26.8521
R2223 VDD.n2987 VDD.n2939 26.8521
R2224 VDD.n2987 VDD.n2937 26.8521
R2225 VDD.n2987 VDD.n2934 26.8521
R2226 VDD.n2987 VDD.n2931 26.8521
R2227 VDD.n2987 VDD.n2928 26.8521
R2228 VDD.n2987 VDD.n2925 26.8521
R2229 VDD.n2987 VDD.n2922 26.8521
R2230 VDD.n2987 VDD.n2919 26.8521
R2231 VDD.n2987 VDD.n2916 26.8521
R2232 VDD.n2987 VDD.n2913 26.8521
R2233 VDD.n2987 VDD.n2910 26.8521
R2234 VDD.n2987 VDD.n2907 26.8521
R2235 VDD.n2987 VDD.n2904 26.8521
R2236 VDD.n2987 VDD.n2901 26.8521
R2237 VDD.n2987 VDD.n2900 26.8521
R2238 VDD.n2987 VDD.n2899 26.8521
R2239 VDD.n1232 VDD.n1231 26.8521
R2240 VDD.n1231 VDD.n1230 26.8521
R2241 VDD.n5261 VDD.n5233 26.8521
R2242 VDD.n5261 VDD.n5232 26.8521
R2243 VDD.n1252 VDD.n1246 25.6005
R2244 VDD.n1246 VDD.n1244 25.6005
R2245 VDD.n1244 VDD.n1241 25.6005
R2246 VDD.n1241 VDD.n1239 25.6005
R2247 VDD.n1239 VDD.n1237 25.6005
R2248 VDD.n1709 VDD.n1703 25.6005
R2249 VDD.n1703 VDD.n1701 25.6005
R2250 VDD.n1701 VDD.n1698 25.6005
R2251 VDD.n1698 VDD.n1696 25.6005
R2252 VDD.n1696 VDD.n1694 25.6005
R2253 VDD.n1687 VDD.n1681 25.6005
R2254 VDD.n1681 VDD.n1679 25.6005
R2255 VDD.n1679 VDD.n1676 25.6005
R2256 VDD.n1676 VDD.n1674 25.6005
R2257 VDD.n1674 VDD.n1672 25.6005
R2258 VDD.n1553 VDD.n1547 25.6005
R2259 VDD.n1547 VDD.n1545 25.6005
R2260 VDD.n1545 VDD.n1542 25.6005
R2261 VDD.n1542 VDD.n1540 25.6005
R2262 VDD.n1540 VDD.n1538 25.6005
R2263 VDD.n1571 VDD.n1565 25.6005
R2264 VDD.n1565 VDD.n1563 25.6005
R2265 VDD.n1563 VDD.n1560 25.6005
R2266 VDD.n1560 VDD.n1558 25.6005
R2267 VDD.n1558 VDD.n1556 25.6005
R2268 VDD.n1234 VDD.n1228 25.6005
R2269 VDD.n1228 VDD.n1226 25.6005
R2270 VDD.n1226 VDD.n1223 25.6005
R2271 VDD.n1325 VDD.n1322 25.6005
R2272 VDD.n1445 VDD.n1439 25.6005
R2273 VDD.n1439 VDD.n1436 25.6005
R2274 VDD.n1436 VDD.n1433 25.6005
R2275 VDD.n1433 VDD.n1430 25.6005
R2276 VDD.n3482 VDD.n3475 25.5522
R2277 VDD.n3572 VDD.n3565 25.5522
R2278 VDD.n3846 VDD.n3839 25.5522
R2279 VDD.n3931 VDD.n3924 25.5522
R2280 VDD.n4192 VDD.n4187 25.5522
R2281 VDD.n4264 VDD.n4259 25.5522
R2282 VDD.n4523 VDD.n4514 25.5522
R2283 VDD.n4598 VDD.n4591 25.5522
R2284 VDD.n4873 VDD.n4866 25.5522
R2285 VDD.n4956 VDD.n4949 25.5522
R2286 VDD.n881 VDD.n880 25.3507
R2287 VDD.n6494 VDD.n6493 25.3507
R2288 VDD.n6500 VDD.n6499 25.3505
R2289 VDD.n867 VDD.n866 25.3505
R2290 VDD.n3393 VDD.n3392 23.5867
R2291 VDD.n3648 VDD.n3647 23.5867
R2292 VDD.n3755 VDD.n3754 23.5867
R2293 VDD.n4012 VDD.n4011 23.5867
R2294 VDD.n4109 VDD.n4108 23.5867
R2295 VDD.n4339 VDD.n4338 23.5867
R2296 VDD.n4430 VDD.n4429 23.5867
R2297 VDD.n4683 VDD.n4682 23.5867
R2298 VDD.n4777 VDD.n4776 23.5867
R2299 VDD.n5036 VDD.n5035 23.5867
R2300 VDD.n5132 VDD.n5131 23.5867
R2301 VDD.n3461 VDD.n3454 21.6212
R2302 VDD.n3592 VDD.n3585 21.6212
R2303 VDD.n3823 VDD.n3816 21.6212
R2304 VDD.n3952 VDD.n3945 21.6212
R2305 VDD.n4173 VDD.n4167 21.6212
R2306 VDD.n4280 VDD.n4275 21.6212
R2307 VDD.n4499 VDD.n4492 21.6212
R2308 VDD.n4622 VDD.n4615 21.6212
R2309 VDD.n4854 VDD.n4849 21.6212
R2310 VDD.n4979 VDD.n4972 21.6212
R2311 VDD.n1414 VDD.n1412 19.8574
R2312 VDD.n3413 VDD.n3412 19.6557
R2313 VDD.n3624 VDD.n3623 19.6557
R2314 VDD.n3775 VDD.n3774 19.6557
R2315 VDD.n3988 VDD.n3987 19.6557
R2316 VDD.n4127 VDD.n4126 19.6557
R2317 VDD.n4318 VDD.n4317 19.6557
R2318 VDD.n4448 VDD.n4447 19.6557
R2319 VDD.n4661 VDD.n4660 19.6557
R2320 VDD.n4800 VDD.n4799 19.6557
R2321 VDD.n5017 VDD.n5016 19.6557
R2322 VDD.n5154 VDD.n5153 19.6557
R2323 VDD.n1357 VDD.n1355 18.4588
R2324 VDD.n3441 VDD.n3434 17.6902
R2325 VDD.n3613 VDD.n3606 17.6902
R2326 VDD.n3802 VDD.n3795 17.6902
R2327 VDD.n3970 VDD.n3963 17.6902
R2328 VDD.n4151 VDD.n4146 17.6902
R2329 VDD.n4301 VDD.n4296 17.6902
R2330 VDD.n4475 VDD.n4468 17.6902
R2331 VDD.n4645 VDD.n4638 17.6902
R2332 VDD.n4833 VDD.n4824 17.6902
R2333 VDD.n5003 VDD.n4996 17.6902
R2334 VDD.n1347 VDD.n1346 17.1609
R2335 VDD.n1336 VDD.n1334 17.1609
R2336 VDD.n1334 VDD.n1333 17.1609
R2337 VDD.n1691 VDD.n1688 17.1609
R2338 VDD.n1691 VDD.n1690 17.1609
R2339 VDD.n1669 VDD.n1665 17.1609
R2340 VDD.n1669 VDD.n1668 17.1609
R2341 VDD.n1535 VDD.n1532 17.1609
R2342 VDD.n1535 VDD.n1534 17.1609
R2343 VDD.n1387 VDD.n1386 17.1609
R2344 VDD.n1389 VDD.n1387 17.1609
R2345 VDD.n1400 VDD.n1399 17.1609
R2346 VDD.n1402 VDD.n1400 17.1609
R2347 VDD.n3434 VDD.n3433 15.7246
R2348 VDD.n3606 VDD.n3605 15.7246
R2349 VDD.n3795 VDD.n3794 15.7246
R2350 VDD.n3963 VDD.n3962 15.7246
R2351 VDD.n4146 VDD.n4145 15.7246
R2352 VDD.n4296 VDD.n4295 15.7246
R2353 VDD.n4468 VDD.n4467 15.7246
R2354 VDD.n4638 VDD.n4637 15.7246
R2355 VDD.n4824 VDD.n4823 15.7246
R2356 VDD.n4996 VDD.n4995 15.7246
R2357 VDD.n1349 VDD.n1347 15.6137
R2358 VDD.n3420 VDD.n3413 13.7591
R2359 VDD.n3631 VDD.n3624 13.7591
R2360 VDD.n3782 VDD.n3775 13.7591
R2361 VDD.n3995 VDD.n3988 13.7591
R2362 VDD.n4132 VDD.n4127 13.7591
R2363 VDD.n4323 VDD.n4318 13.7591
R2364 VDD.n4454 VDD.n4448 13.7591
R2365 VDD.n4668 VDD.n4661 13.7591
R2366 VDD.n4807 VDD.n4800 13.7591
R2367 VDD.n5024 VDD.n5017 13.7591
R2368 VDD.n5264 VDD.n5154 13.7591
R2369 VDD.n103 VDD.n102 13.177
R2370 VDD.n2289 VDD.n2288 13.1521
R2371 VDD.n2282 VDD.n2281 13.1521
R2372 VDD.n2275 VDD.n2274 13.1521
R2373 VDD.n2268 VDD.n2267 13.1521
R2374 VDD.n2261 VDD.n2260 13.1521
R2375 VDD.n2254 VDD.n2253 13.1521
R2376 VDD.n2247 VDD.n2246 13.1521
R2377 VDD.n2240 VDD.n2239 13.1521
R2378 VDD.n2233 VDD.n2232 13.1521
R2379 VDD.n2226 VDD.n2225 13.1521
R2380 VDD.n2219 VDD.n2218 13.1521
R2381 VDD.n2212 VDD.n2211 13.1521
R2382 VDD.n2205 VDD.n2204 13.1521
R2383 VDD.n2198 VDD.n2197 13.1521
R2384 VDD.n2191 VDD.n2190 13.1521
R2385 VDD.n2184 VDD.n2183 13.1521
R2386 VDD.n2177 VDD.n2176 13.1521
R2387 VDD.n2170 VDD.n2169 13.1521
R2388 VDD.n2163 VDD.n2162 13.1521
R2389 VDD.n2156 VDD.n2155 13.1521
R2390 VDD.n2647 VDD.n2646 13.1515
R2391 VDD.n2640 VDD.n2639 13.1515
R2392 VDD.n2633 VDD.n2632 13.1515
R2393 VDD.n2626 VDD.n2625 13.1515
R2394 VDD.n2619 VDD.n2618 13.1515
R2395 VDD.n2612 VDD.n2611 13.1515
R2396 VDD.n2605 VDD.n2604 13.1515
R2397 VDD.n2598 VDD.n2597 13.1515
R2398 VDD.n2591 VDD.n2590 13.1515
R2399 VDD.n2584 VDD.n2583 13.1515
R2400 VDD.n2577 VDD.n2576 13.1515
R2401 VDD.n2570 VDD.n2569 13.1515
R2402 VDD.n2563 VDD.n2562 13.1515
R2403 VDD.n2556 VDD.n2555 13.1515
R2404 VDD.n2549 VDD.n2548 13.1515
R2405 VDD.n2542 VDD.n2541 13.1515
R2406 VDD.n2535 VDD.n2534 13.1515
R2407 VDD.n2528 VDD.n2527 13.1515
R2408 VDD.n2521 VDD.n2520 13.1515
R2409 VDD.n2514 VDD.n2513 13.1515
R2410 VDD.n2468 VDD.n2467 13.1515
R2411 VDD.n2461 VDD.n2460 13.1515
R2412 VDD.n2454 VDD.n2453 13.1515
R2413 VDD.n2447 VDD.n2446 13.1515
R2414 VDD.n2440 VDD.n2439 13.1515
R2415 VDD.n2433 VDD.n2432 13.1515
R2416 VDD.n2426 VDD.n2425 13.1515
R2417 VDD.n2419 VDD.n2418 13.1515
R2418 VDD.n2412 VDD.n2411 13.1515
R2419 VDD.n2405 VDD.n2404 13.1515
R2420 VDD.n2398 VDD.n2397 13.1515
R2421 VDD.n2391 VDD.n2390 13.1515
R2422 VDD.n2384 VDD.n2383 13.1515
R2423 VDD.n2377 VDD.n2376 13.1515
R2424 VDD.n2370 VDD.n2369 13.1515
R2425 VDD.n2363 VDD.n2362 13.1515
R2426 VDD.n2356 VDD.n2355 13.1515
R2427 VDD.n2349 VDD.n2348 13.1515
R2428 VDD.n2342 VDD.n2341 13.1515
R2429 VDD.n2335 VDD.n2334 13.1515
R2430 VDD.n2113 VDD.n2112 13.1509
R2431 VDD.n2106 VDD.n2105 13.1509
R2432 VDD.n2099 VDD.n2098 13.1509
R2433 VDD.n2092 VDD.n2091 13.1509
R2434 VDD.n2085 VDD.n2084 13.1509
R2435 VDD.n2078 VDD.n2077 13.1509
R2436 VDD.n2071 VDD.n2070 13.1509
R2437 VDD.n2064 VDD.n2063 13.1509
R2438 VDD.n2057 VDD.n2056 13.1509
R2439 VDD.n2050 VDD.n2049 13.1509
R2440 VDD.n2043 VDD.n2042 13.1509
R2441 VDD.n2036 VDD.n2035 13.1509
R2442 VDD.n2029 VDD.n2028 13.1509
R2443 VDD.n2022 VDD.n2021 13.1509
R2444 VDD.n2015 VDD.n2014 13.1509
R2445 VDD.n2008 VDD.n2007 13.1509
R2446 VDD.n2001 VDD.n2000 13.1509
R2447 VDD.n1994 VDD.n1993 13.1509
R2448 VDD.n1987 VDD.n1986 13.1509
R2449 VDD.n1980 VDD.n1979 13.1509
R2450 VDD.n5853 VDD.n5852 13.1501
R2451 VDD.n5846 VDD.n5845 13.1501
R2452 VDD.n5839 VDD.n5838 13.1501
R2453 VDD.n5832 VDD.n5831 13.1501
R2454 VDD.n5825 VDD.n5824 13.1501
R2455 VDD.n5818 VDD.n5817 13.1501
R2456 VDD.n5811 VDD.n5810 13.1501
R2457 VDD.n5804 VDD.n5803 13.1501
R2458 VDD.n5797 VDD.n5796 13.1501
R2459 VDD.n5790 VDD.n5789 13.1501
R2460 VDD.n5783 VDD.n5782 13.1501
R2461 VDD.n5776 VDD.n5775 13.1501
R2462 VDD.n5769 VDD.n5768 13.1501
R2463 VDD.n5762 VDD.n5761 13.1501
R2464 VDD.n5755 VDD.n5754 13.1501
R2465 VDD.n5748 VDD.n5747 13.1501
R2466 VDD.n5741 VDD.n5740 13.1501
R2467 VDD.n5734 VDD.n5733 13.1501
R2468 VDD.n5727 VDD.n5726 13.1501
R2469 VDD.n5720 VDD.n5719 13.1501
R2470 VDD.n1934 VDD.n1933 13.1501
R2471 VDD.n1927 VDD.n1926 13.1501
R2472 VDD.n1920 VDD.n1919 13.1501
R2473 VDD.n1913 VDD.n1912 13.1501
R2474 VDD.n1906 VDD.n1905 13.1501
R2475 VDD.n1899 VDD.n1898 13.1501
R2476 VDD.n1892 VDD.n1891 13.1501
R2477 VDD.n1885 VDD.n1884 13.1501
R2478 VDD.n1878 VDD.n1877 13.1501
R2479 VDD.n1871 VDD.n1870 13.1501
R2480 VDD.n1864 VDD.n1863 13.1501
R2481 VDD.n1857 VDD.n1856 13.1501
R2482 VDD.n1850 VDD.n1849 13.1501
R2483 VDD.n1843 VDD.n1842 13.1501
R2484 VDD.n1836 VDD.n1835 13.1501
R2485 VDD.n1829 VDD.n1828 13.1501
R2486 VDD.n1822 VDD.n1821 13.1501
R2487 VDD.n1815 VDD.n1814 13.1501
R2488 VDD.n1808 VDD.n1807 13.1501
R2489 VDD.n1801 VDD.n1800 13.1501
R2490 VDD.n5674 VDD.n5673 13.1489
R2491 VDD.n5667 VDD.n5666 13.1489
R2492 VDD.n5660 VDD.n5659 13.1489
R2493 VDD.n5653 VDD.n5652 13.1489
R2494 VDD.n5646 VDD.n5645 13.1489
R2495 VDD.n5639 VDD.n5638 13.1489
R2496 VDD.n5632 VDD.n5631 13.1489
R2497 VDD.n5625 VDD.n5624 13.1489
R2498 VDD.n5618 VDD.n5617 13.1489
R2499 VDD.n5611 VDD.n5610 13.1489
R2500 VDD.n5604 VDD.n5603 13.1489
R2501 VDD.n5597 VDD.n5596 13.1489
R2502 VDD.n5590 VDD.n5589 13.1489
R2503 VDD.n5583 VDD.n5582 13.1489
R2504 VDD.n5576 VDD.n5575 13.1489
R2505 VDD.n5569 VDD.n5568 13.1489
R2506 VDD.n5562 VDD.n5561 13.1489
R2507 VDD.n5555 VDD.n5554 13.1489
R2508 VDD.n5548 VDD.n5547 13.1489
R2509 VDD.n5541 VDD.n5540 13.1489
R2510 VDD.n6032 VDD.n6031 13.1451
R2511 VDD.n6025 VDD.n6024 13.1451
R2512 VDD.n6018 VDD.n6017 13.1451
R2513 VDD.n6011 VDD.n6010 13.1451
R2514 VDD.n6004 VDD.n6003 13.1451
R2515 VDD.n5997 VDD.n5996 13.1451
R2516 VDD.n5990 VDD.n5989 13.1451
R2517 VDD.n5983 VDD.n5982 13.1451
R2518 VDD.n5976 VDD.n5975 13.1451
R2519 VDD.n5969 VDD.n5968 13.1451
R2520 VDD.n5962 VDD.n5961 13.1451
R2521 VDD.n5955 VDD.n5954 13.1451
R2522 VDD.n5948 VDD.n5947 13.1451
R2523 VDD.n5941 VDD.n5940 13.1451
R2524 VDD.n5934 VDD.n5933 13.1451
R2525 VDD.n5927 VDD.n5926 13.1451
R2526 VDD.n5920 VDD.n5919 13.1451
R2527 VDD.n5913 VDD.n5912 13.1451
R2528 VDD.n5906 VDD.n5905 13.1451
R2529 VDD.n5899 VDD.n5898 13.1451
R2530 VDD.n6211 VDD.n6210 13.1389
R2531 VDD.n6204 VDD.n6203 13.1389
R2532 VDD.n6197 VDD.n6196 13.1389
R2533 VDD.n6190 VDD.n6189 13.1389
R2534 VDD.n6183 VDD.n6182 13.1389
R2535 VDD.n6176 VDD.n6175 13.1389
R2536 VDD.n6169 VDD.n6168 13.1389
R2537 VDD.n6162 VDD.n6161 13.1389
R2538 VDD.n6155 VDD.n6154 13.1389
R2539 VDD.n6148 VDD.n6147 13.1389
R2540 VDD.n6141 VDD.n6140 13.1389
R2541 VDD.n6134 VDD.n6133 13.1389
R2542 VDD.n6127 VDD.n6126 13.1389
R2543 VDD.n6120 VDD.n6119 13.1389
R2544 VDD.n6113 VDD.n6112 13.1389
R2545 VDD.n6106 VDD.n6105 13.1389
R2546 VDD.n6099 VDD.n6098 13.1389
R2547 VDD.n6092 VDD.n6091 13.1389
R2548 VDD.n6085 VDD.n6084 13.1389
R2549 VDD.n6078 VDD.n6077 13.1389
R2550 VDD.n5495 VDD.n5494 13.1304
R2551 VDD.n5488 VDD.n5487 13.1304
R2552 VDD.n5481 VDD.n5480 13.1304
R2553 VDD.n5474 VDD.n5473 13.1304
R2554 VDD.n5467 VDD.n5466 13.1304
R2555 VDD.n5460 VDD.n5459 13.1304
R2556 VDD.n5453 VDD.n5452 13.1304
R2557 VDD.n5446 VDD.n5445 13.1304
R2558 VDD.n5439 VDD.n5438 13.1304
R2559 VDD.n5432 VDD.n5431 13.1304
R2560 VDD.n5425 VDD.n5424 13.1304
R2561 VDD.n5418 VDD.n5417 13.1304
R2562 VDD.n5411 VDD.n5410 13.1304
R2563 VDD.n5404 VDD.n5403 13.1304
R2564 VDD.n5397 VDD.n5396 13.1304
R2565 VDD.n5390 VDD.n5389 13.1304
R2566 VDD.n5383 VDD.n5382 13.1304
R2567 VDD.n5376 VDD.n5375 13.1304
R2568 VDD.n5369 VDD.n5368 13.1304
R2569 VDD.n5362 VDD.n5361 13.1304
R2570 VDD.n2896 VDD.n2894 12.4836
R2571 VDD.n2898 VDD.n2896 12.4836
R2572 VDD.n2991 VDD.n2989 12.4836
R2573 VDD.n5200 VDD.n5199 12.4836
R2574 VDD.n5199 VDD.n5198 12.4836
R2575 VDD.n5198 VDD.n5197 12.4836
R2576 VDD.n3454 VDD.n3453 11.7936
R2577 VDD.n3585 VDD.n3584 11.7936
R2578 VDD.n3816 VDD.n3815 11.7936
R2579 VDD.n3945 VDD.n3944 11.7936
R2580 VDD.n4167 VDD.n4166 11.7936
R2581 VDD.n4275 VDD.n4274 11.7936
R2582 VDD.n4492 VDD.n4491 11.7936
R2583 VDD.n4615 VDD.n4614 11.7936
R2584 VDD.n4849 VDD.n4848 11.7936
R2585 VDD.n4972 VDD.n4971 11.7936
R2586 VDD.n4527 VDD.n4526 11.5205
R2587 VDD.n4228 VDD.n4225 10.8805
R2588 VDD.n4228 VDD.n4227 10.8805
R2589 VDD.n4556 VDD.n4553 10.8805
R2590 VDD.n4556 VDD.n4555 10.8805
R2591 VDD.n4911 VDD.n4908 10.8805
R2592 VDD.n4911 VDD.n4910 10.8805
R2593 VDD.n2987 VDD.n2898 10.2807
R2594 VDD.n142 VDD.n141 10.2648
R2595 VDD.n150 VDD.n144 10.2648
R2596 VDD.n148 VDD.n145 10.2648
R2597 VDD.n152 VDD.n143 10.2568
R2598 VDD.n147 VDD.n146 10.1884
R2599 VDD.n2892 VDD.n2891 10.0971
R2600 VDD.n5196 VDD.n5195 9.91354
R2601 VDD.n3400 VDD.n3393 9.82809
R2602 VDD.n3655 VDD.n3648 9.82809
R2603 VDD.n3762 VDD.n3755 9.82809
R2604 VDD.n4019 VDD.n4012 9.82809
R2605 VDD.n4114 VDD.n4109 9.82809
R2606 VDD.n4344 VDD.n4339 9.82809
R2607 VDD.n4435 VDD.n4430 9.82809
R2608 VDD.n4690 VDD.n4683 9.82809
R2609 VDD.n4784 VDD.n4777 9.82809
R2610 VDD.n5043 VDD.n5036 9.82809
R2611 VDD.n5137 VDD.n5132 9.82809
R2612 VDD.n3883 VDD.n3882 9.6005
R2613 VDD.n3893 VDD.n3892 9.6005
R2614 VDD.n1355 VDD.n1353 9.56533
R2615 VDD.n1353 VDD.n1351 9.56533
R2616 VDD.n1351 VDD.n1349 9.56533
R2617 VDD.n1346 VDD.n1344 9.56533
R2618 VDD.n1344 VDD.n1342 9.56533
R2619 VDD.n1342 VDD.n1340 9.56533
R2620 VDD.n1340 VDD.n1338 9.56533
R2621 VDD.n1338 VDD.n1336 9.56533
R2622 VDD.n1333 VDD.n1331 9.56533
R2623 VDD.n1331 VDD.n1329 9.56533
R2624 VDD.n1329 VDD.n1327 9.56533
R2625 VDD.n1327 VDD.n1326 9.56533
R2626 VDD.n1690 VDD.n1689 9.56533
R2627 VDD.n1663 VDD.n1662 9.56533
R2628 VDD.n1664 VDD.n1663 9.56533
R2629 VDD.n1665 VDD.n1664 9.56533
R2630 VDD.n1668 VDD.n1667 9.56533
R2631 VDD.n1667 VDD.n1666 9.56533
R2632 VDD.n1531 VDD.n1530 9.56533
R2633 VDD.n1532 VDD.n1531 9.56533
R2634 VDD.n1534 VDD.n1533 9.56533
R2635 VDD.n1383 VDD.n1382 9.56533
R2636 VDD.n1384 VDD.n1383 9.56533
R2637 VDD.n1386 VDD.n1384 9.56533
R2638 VDD.n1391 VDD.n1389 9.56533
R2639 VDD.n1393 VDD.n1391 9.56533
R2640 VDD.n1395 VDD.n1393 9.56533
R2641 VDD.n1397 VDD.n1395 9.56533
R2642 VDD.n1399 VDD.n1397 9.56533
R2643 VDD.n1404 VDD.n1402 9.56533
R2644 VDD.n1406 VDD.n1404 9.56533
R2645 VDD.n1408 VDD.n1406 9.56533
R2646 VDD.n1410 VDD.n1408 9.56533
R2647 VDD.n1412 VDD.n1410 9.56533
R2648 VDD.n108 VDD.n107 9.3182
R2649 VDD.n4050 VDD.n4049 9.3005
R2650 VDD.n4083 VDD.n4082 9.3005
R2651 VDD.n4353 VDD.n4352 9.3005
R2652 VDD.n4372 VDD.n4371 9.3005
R2653 VDD.n4404 VDD.n4403 9.3005
R2654 VDD.n4440 VDD.n4439 9.3005
R2655 VDD.n4679 VDD.n4678 9.3005
R2656 VDD.n4718 VDD.n4717 9.3005
R2657 VDD.n4753 VDD.n4752 9.3005
R2658 VDD.n5072 VDD.n5071 9.3005
R2659 VDD.n5106 VDD.n5105 9.3005
R2660 VDD.n5011 VDD.n5010 9.3005
R2661 VDD.n4921 VDD.n4920 9.3005
R2662 VDD.n4846 VDD.n4845 9.3005
R2663 VDD.n4677 VDD.n4676 9.3005
R2664 VDD.n4604 VDD.n4603 9.3005
R2665 VDD.n4442 VDD.n4441 9.3005
R2666 VDD.n4355 VDD.n4354 9.3005
R2667 VDD.n4288 VDD.n4287 9.3005
R2668 VDD.n4217 VDD.n4216 9.3005
R2669 VDD.n4139 VDD.n4138 9.3005
R2670 VDD.n4052 VDD.n4051 9.3005
R2671 VDD.n3978 VDD.n3977 9.3005
R2672 VDD.n3888 VDD.n3887 9.3005
R2673 VDD.n3809 VDD.n3808 9.3005
R2674 VDD.n3712 VDD.n3711 9.3005
R2675 VDD.n3638 VDD.n3637 9.3005
R2676 VDD.n3536 VDD.n3535 9.3005
R2677 VDD.n3468 VDD.n3467 9.3005
R2678 VDD.n3023 VDD.n3022 9.3005
R2679 VDD.n5104 VDD.n5103 9.3005
R2680 VDD.n2997 VDD.n2996 9.3005
R2681 VDD.n2996 VDD.n2995 9.3005
R2682 VDD.n3037 VDD.n3036 9.3005
R2683 VDD.n3036 VDD.n3035 9.3005
R2684 VDD.n3016 VDD.n3015 9.3005
R2685 VDD.n3015 VDD.n3014 9.3005
R2686 VDD.n3401 VDD.n3400 9.3005
R2687 VDD.n3400 VDD.n3399 9.3005
R2688 VDD.n3421 VDD.n3420 9.3005
R2689 VDD.n3420 VDD.n3419 9.3005
R2690 VDD.n3442 VDD.n3441 9.3005
R2691 VDD.n3441 VDD.n3440 9.3005
R2692 VDD.n3462 VDD.n3461 9.3005
R2693 VDD.n3461 VDD.n3460 9.3005
R2694 VDD.n3483 VDD.n3482 9.3005
R2695 VDD.n3482 VDD.n3481 9.3005
R2696 VDD.n3510 VDD.n3509 9.3005
R2697 VDD.n3509 VDD.n3508 9.3005
R2698 VDD.n3554 VDD.n3553 9.3005
R2699 VDD.n3553 VDD.n3552 9.3005
R2700 VDD.n3573 VDD.n3572 9.3005
R2701 VDD.n3572 VDD.n3571 9.3005
R2702 VDD.n3593 VDD.n3592 9.3005
R2703 VDD.n3592 VDD.n3591 9.3005
R2704 VDD.n3614 VDD.n3613 9.3005
R2705 VDD.n3613 VDD.n3612 9.3005
R2706 VDD.n3632 VDD.n3631 9.3005
R2707 VDD.n3631 VDD.n3630 9.3005
R2708 VDD.n3656 VDD.n3655 9.3005
R2709 VDD.n3655 VDD.n3654 9.3005
R2710 VDD.n3680 VDD.n3679 9.3005
R2711 VDD.n3679 VDD.n3678 9.3005
R2712 VDD.n3703 VDD.n3702 9.3005
R2713 VDD.n3702 VDD.n3701 9.3005
R2714 VDD.n3724 VDD.n3723 9.3005
R2715 VDD.n3723 VDD.n3722 9.3005
R2716 VDD.n3743 VDD.n3742 9.3005
R2717 VDD.n3742 VDD.n3741 9.3005
R2718 VDD.n3763 VDD.n3762 9.3005
R2719 VDD.n3762 VDD.n3761 9.3005
R2720 VDD.n3783 VDD.n3782 9.3005
R2721 VDD.n3782 VDD.n3781 9.3005
R2722 VDD.n3803 VDD.n3802 9.3005
R2723 VDD.n3802 VDD.n3801 9.3005
R2724 VDD.n3824 VDD.n3823 9.3005
R2725 VDD.n3823 VDD.n3822 9.3005
R2726 VDD.n3847 VDD.n3846 9.3005
R2727 VDD.n3846 VDD.n3845 9.3005
R2728 VDD.n3876 VDD.n3875 9.3005
R2729 VDD.n3875 VDD.n3874 9.3005
R2730 VDD.n3916 VDD.n3915 9.3005
R2731 VDD.n3915 VDD.n3914 9.3005
R2732 VDD.n3914 VDD.n3913 9.3005
R2733 VDD.n3932 VDD.n3931 9.3005
R2734 VDD.n3931 VDD.n3930 9.3005
R2735 VDD.n3953 VDD.n3952 9.3005
R2736 VDD.n3952 VDD.n3951 9.3005
R2737 VDD.n3971 VDD.n3970 9.3005
R2738 VDD.n3970 VDD.n3969 9.3005
R2739 VDD.n3996 VDD.n3995 9.3005
R2740 VDD.n3995 VDD.n3994 9.3005
R2741 VDD.n4020 VDD.n4019 9.3005
R2742 VDD.n4019 VDD.n4018 9.3005
R2743 VDD.n4042 VDD.n4041 9.3005
R2744 VDD.n4041 VDD.n4040 9.3005
R2745 VDD.n4061 VDD.n4060 9.3005
R2746 VDD.n4060 VDD.n4059 9.3005
R2747 VDD.n4078 VDD.n4077 9.3005
R2748 VDD.n4077 VDD.n4076 9.3005
R2749 VDD.n4096 VDD.n4095 9.3005
R2750 VDD.n4095 VDD.n4094 9.3005
R2751 VDD.n4115 VDD.n4114 9.3005
R2752 VDD.n4114 VDD.n4113 9.3005
R2753 VDD.n4133 VDD.n4132 9.3005
R2754 VDD.n4132 VDD.n4131 9.3005
R2755 VDD.n4152 VDD.n4151 9.3005
R2756 VDD.n4151 VDD.n4150 9.3005
R2757 VDD.n4174 VDD.n4173 9.3005
R2758 VDD.n4173 VDD.n4172 9.3005
R2759 VDD.n4193 VDD.n4192 9.3005
R2760 VDD.n4192 VDD.n4191 9.3005
R2761 VDD.n4215 VDD.n4214 9.3005
R2762 VDD.n4214 VDD.n4213 9.3005
R2763 VDD.n4213 VDD.n4212 9.3005
R2764 VDD.n4250 VDD.n4249 9.3005
R2765 VDD.n4249 VDD.n4248 9.3005
R2766 VDD.n4248 VDD.n4247 9.3005
R2767 VDD.n4265 VDD.n4264 9.3005
R2768 VDD.n4264 VDD.n4263 9.3005
R2769 VDD.n4281 VDD.n4280 9.3005
R2770 VDD.n4280 VDD.n4279 9.3005
R2771 VDD.n4302 VDD.n4301 9.3005
R2772 VDD.n4301 VDD.n4300 9.3005
R2773 VDD.n4324 VDD.n4323 9.3005
R2774 VDD.n4323 VDD.n4322 9.3005
R2775 VDD.n4345 VDD.n4344 9.3005
R2776 VDD.n4344 VDD.n4343 9.3005
R2777 VDD.n4364 VDD.n4363 9.3005
R2778 VDD.n4363 VDD.n4362 9.3005
R2779 VDD.n4382 VDD.n4381 9.3005
R2780 VDD.n4381 VDD.n4380 9.3005
R2781 VDD.n4399 VDD.n4398 9.3005
R2782 VDD.n4398 VDD.n4397 9.3005
R2783 VDD.n4418 VDD.n4417 9.3005
R2784 VDD.n4417 VDD.n4416 9.3005
R2785 VDD.n4436 VDD.n4435 9.3005
R2786 VDD.n4435 VDD.n4434 9.3005
R2787 VDD.n4455 VDD.n4454 9.3005
R2788 VDD.n4454 VDD.n4453 9.3005
R2789 VDD.n4476 VDD.n4475 9.3005
R2790 VDD.n4475 VDD.n4474 9.3005
R2791 VDD.n4500 VDD.n4499 9.3005
R2792 VDD.n4499 VDD.n4498 9.3005
R2793 VDD.n4524 VDD.n4523 9.3005
R2794 VDD.n4523 VDD.n4522 9.3005
R2795 VDD.n4544 VDD.n4543 9.3005
R2796 VDD.n4543 VDD.n4542 9.3005
R2797 VDD.n4582 VDD.n4581 9.3005
R2798 VDD.n4581 VDD.n4580 9.3005
R2799 VDD.n4580 VDD.n4579 9.3005
R2800 VDD.n4600 VDD.n4599 9.3005
R2801 VDD.n4599 VDD.n4598 9.3005
R2802 VDD.n4598 VDD.n4597 9.3005
R2803 VDD.n4623 VDD.n4622 9.3005
R2804 VDD.n4622 VDD.n4621 9.3005
R2805 VDD.n4646 VDD.n4645 9.3005
R2806 VDD.n4645 VDD.n4644 9.3005
R2807 VDD.n4669 VDD.n4668 9.3005
R2808 VDD.n4668 VDD.n4667 9.3005
R2809 VDD.n4691 VDD.n4690 9.3005
R2810 VDD.n4690 VDD.n4689 9.3005
R2811 VDD.n4710 VDD.n4709 9.3005
R2812 VDD.n4709 VDD.n4708 9.3005
R2813 VDD.n4730 VDD.n4729 9.3005
R2814 VDD.n4729 VDD.n4728 9.3005
R2815 VDD.n4749 VDD.n4748 9.3005
R2816 VDD.n4748 VDD.n4747 9.3005
R2817 VDD.n4768 VDD.n4767 9.3005
R2818 VDD.n4767 VDD.n4766 9.3005
R2819 VDD.n4785 VDD.n4784 9.3005
R2820 VDD.n4784 VDD.n4783 9.3005
R2821 VDD.n4808 VDD.n4807 9.3005
R2822 VDD.n4807 VDD.n4806 9.3005
R2823 VDD.n4834 VDD.n4833 9.3005
R2824 VDD.n4833 VDD.n4832 9.3005
R2825 VDD.n4855 VDD.n4854 9.3005
R2826 VDD.n4854 VDD.n4853 9.3005
R2827 VDD.n4874 VDD.n4873 9.3005
R2828 VDD.n4873 VDD.n4872 9.3005
R2829 VDD.n4898 VDD.n4897 9.3005
R2830 VDD.n4897 VDD.n4896 9.3005
R2831 VDD.n4938 VDD.n4937 9.3005
R2832 VDD.n4937 VDD.n4936 9.3005
R2833 VDD.n4936 VDD.n4935 9.3005
R2834 VDD.n4957 VDD.n4956 9.3005
R2835 VDD.n4956 VDD.n4955 9.3005
R2836 VDD.n4980 VDD.n4979 9.3005
R2837 VDD.n4979 VDD.n4978 9.3005
R2838 VDD.n5004 VDD.n5003 9.3005
R2839 VDD.n5003 VDD.n5002 9.3005
R2840 VDD.n5025 VDD.n5024 9.3005
R2841 VDD.n5024 VDD.n5023 9.3005
R2842 VDD.n5044 VDD.n5043 9.3005
R2843 VDD.n5043 VDD.n5042 9.3005
R2844 VDD.n5064 VDD.n5063 9.3005
R2845 VDD.n5063 VDD.n5062 9.3005
R2846 VDD.n5083 VDD.n5082 9.3005
R2847 VDD.n5082 VDD.t120 9.3005
R2848 VDD.n5098 VDD.n5097 9.3005
R2849 VDD.n5097 VDD.n5096 9.3005
R2850 VDD.n5117 VDD.n5116 9.3005
R2851 VDD.n5116 VDD.n5115 9.3005
R2852 VDD.n5138 VDD.n5137 9.3005
R2853 VDD.n5137 VDD.n5136 9.3005
R2854 VDD.n5265 VDD.n5264 9.3005
R2855 VDD.n5264 VDD.n5263 9.3005
R2856 VDD.n92 VDD.n91 9.3005
R2857 VDD.n3548 VDD.n3546 9.17924
R2858 VDD.n3909 VDD.n3907 9.17924
R2859 VDD.n4244 VDD.n4243 9.17924
R2860 VDD.n4931 VDD.n4929 9.17924
R2861 VDD.n107 VDD.n106 9.0206
R2862 VDD.n5262 VDD.n5261 8.81209
R2863 VDD.n3531 VDD.n3530 8.3205
R2864 VDD.n5263 VDD.n5262 7.89422
R2865 VDD.n3475 VDD.n3474 7.86257
R2866 VDD.n3565 VDD.n3564 7.86257
R2867 VDD.n3839 VDD.n3838 7.86257
R2868 VDD.n3924 VDD.n3923 7.86257
R2869 VDD.n4187 VDD.n4186 7.86257
R2870 VDD.n4259 VDD.n4258 7.86257
R2871 VDD.n4514 VDD.n4513 7.86257
R2872 VDD.n4591 VDD.n4590 7.86257
R2873 VDD.n4866 VDD.n4865 7.86257
R2874 VDD.n4949 VDD.n4948 7.86257
R2875 VDD.n4832 VDD.n4831 7.52707
R2876 VDD.n1526 VDD.n1378 7.44755
R2877 VDD.n1527 VDD.n1377 7.44755
R2878 VDD.n1528 VDD.n1376 7.44755
R2879 VDD.n1529 VDD.n1375 7.44755
R2880 VDD.n1374 VDD.n1209 7.29594
R2881 VDD.n4172 VDD.n4171 7.15992
R2882 VDD.n4522 VDD.n4521 6.79277
R2883 VDD.n3874 VDD.n3873 6.42562
R2884 VDD.n4212 VDD.n4211 6.42562
R2885 VDD.n4542 VDD.n4541 6.42562
R2886 VDD.n3524 VDD.n3522 6.0805
R2887 VDD.t19 VDD.n3869 6.05847
R2888 VDD.n3015 VDD.n3008 5.89705
R2889 VDD.n3679 VDD.n3672 5.89705
R2890 VDD.n3742 VDD.n3735 5.89705
R2891 VDD.n4041 VDD.n4035 5.89705
R2892 VDD.n4095 VDD.n4090 5.89705
R2893 VDD.n4363 VDD.n4358 5.89705
R2894 VDD.n4417 VDD.n4412 5.89705
R2895 VDD.n4709 VDD.n4702 5.89705
R2896 VDD.n4767 VDD.n4760 5.89705
R2897 VDD.n5063 VDD.n5056 5.89705
R2898 VDD.n5116 VDD.n5111 5.89705
R2899 VDD.n4896 VDD.t83 5.8749
R2900 VDD.n2998 VDD.n2833 5.80588
R2901 VDD.n3508 VDD.t45 5.50775
R2902 VDD.t21 VDD.n4573 5.32417
R2903 VDD.n6749 VDD.n6746 5.27565
R2904 VDD.n6746 VDD.n6743 5.27565
R2905 VDD.n6743 VDD.n6740 5.27565
R2906 VDD.n6740 VDD.n6737 5.27565
R2907 VDD.n6737 VDD.n6734 5.27565
R2908 VDD.n6734 VDD.n6731 5.27565
R2909 VDD.n6731 VDD.n6728 5.27565
R2910 VDD.n6728 VDD.n6725 5.27565
R2911 VDD.n6725 VDD.n6722 5.27565
R2912 VDD.n6722 VDD.n6719 5.27565
R2913 VDD.n175 VDD.n172 5.27565
R2914 VDD.n267 VDD.n264 5.27565
R2915 VDD.n270 VDD.n267 5.27565
R2916 VDD.n273 VDD.n270 5.27565
R2917 VDD.n276 VDD.n273 5.27565
R2918 VDD.n279 VDD.n276 5.27565
R2919 VDD.n282 VDD.n279 5.27565
R2920 VDD.n285 VDD.n282 5.27565
R2921 VDD.n288 VDD.n285 5.27565
R2922 VDD.n1207 VDD.n1018 5.19794
R2923 VDD.n4070 VDD.n4069 5.1205
R2924 VDD.n4374 VDD.n4373 5.1205
R2925 VDD.n4391 VDD.n4390 5.1205
R2926 VDD.n4720 VDD.n4719 5.1205
R2927 VDD.n4739 VDD.n4738 5.1205
R2928 VDD.n5075 VDD.n5074 5.1205
R2929 VDD.n1155 VDD.n1152 5.1205
R2930 VDD.n1152 VDD.n1149 5.1205
R2931 VDD.n1149 VDD.n1146 5.1205
R2932 VDD.n1146 VDD.n1143 5.1205
R2933 VDD.n1143 VDD.n1140 5.1205
R2934 VDD.n1140 VDD.n1137 5.1205
R2935 VDD.n1137 VDD.n1134 5.1205
R2936 VDD.n1134 VDD.n1131 5.1205
R2937 VDD.n1131 VDD.n1128 5.1205
R2938 VDD.n1128 VDD.n1125 5.1205
R2939 VDD.n1125 VDD.n1122 5.1205
R2940 VDD.n1122 VDD.n1119 5.1205
R2941 VDD.n1119 VDD.n1116 5.1205
R2942 VDD.n1116 VDD.n1113 5.1205
R2943 VDD.n1113 VDD.n1110 5.1205
R2944 VDD.n1110 VDD.n1107 5.1205
R2945 VDD.n953 VDD.n950 5.1205
R2946 VDD.n956 VDD.n953 5.1205
R2947 VDD.n959 VDD.n956 5.1205
R2948 VDD.n962 VDD.n959 5.1205
R2949 VDD.n965 VDD.n962 5.1205
R2950 VDD.n968 VDD.n965 5.1205
R2951 VDD.n971 VDD.n968 5.1205
R2952 VDD.n974 VDD.n971 5.1205
R2953 VDD.n977 VDD.n974 5.1205
R2954 VDD.n980 VDD.n977 5.1205
R2955 VDD.n983 VDD.n980 5.1205
R2956 VDD.n986 VDD.n983 5.1205
R2957 VDD.n989 VDD.n986 5.1205
R2958 VDD.n992 VDD.n989 5.1205
R2959 VDD.n995 VDD.n992 5.1205
R2960 VDD.n998 VDD.n995 5.1205
R2961 VDD.n1001 VDD.n998 5.1205
R2962 VDD.n1004 VDD.n1001 5.1205
R2963 VDD.n1007 VDD.n1004 5.1205
R2964 VDD.n1010 VDD.n1007 5.1205
R2965 VDD.n1013 VDD.n1010 5.1205
R2966 VDD.n1016 VDD.n1013 5.1205
R2967 VDD.n885 VDD.n882 5.1205
R2968 VDD.n3510 VDD.n3496 4.8005
R2969 VDD.n3554 VDD.n3540 4.8005
R2970 VDD.n3876 VDD.n3859 4.8005
R2971 VDD.n3915 VDD.n3903 4.8005
R2972 VDD.n4214 VDD.n4205 4.8005
R2973 VDD.n4249 VDD.n4239 4.8005
R2974 VDD.n4544 VDD.n4532 4.8005
R2975 VDD.n4546 VDD.n4544 4.8005
R2976 VDD.n4581 VDD.n4567 4.8005
R2977 VDD.n4857 VDD.n4855 4.8005
R2978 VDD.n4898 VDD.n4884 4.8005
R2979 VDD.n4900 VDD.n4898 4.8005
R2980 VDD.n4937 VDD.n4923 4.8005
R2981 VDD.n5100 VDD.n5090 4.8005
R2982 VDD.n4434 VDD.t70 4.77345
R2983 VDD.n292 VDD.n288 4.73262
R2984 VDD.n5354 VDD.n5353 4.72967
R2985 VDD.n6265 VDD.n6259 4.7192
R2986 VDD.n181 VDD.n176 4.71572
R2987 VDD.n261 VDD.n260 4.71572
R2988 VDD.n297 VDD.n292 4.71572
R2989 VDD.n4771 VDD.n4770 4.6505
R2990 VDD.n4303 VDD.n4302 4.6505
R2991 VDD.n4525 VDD.n4524 4.6505
R2992 VDD.n5266 VDD.n5265 4.6505
R2993 VDD.n904 VDD.n903 4.6505
R2994 VDD.n909 VDD.n908 4.6505
R2995 VDD.n914 VDD.n913 4.6505
R2996 VDD.n922 VDD.n921 4.6505
R2997 VDD.n927 VDD.n926 4.6505
R2998 VDD.n932 VDD.n931 4.6505
R2999 VDD.n937 VDD.n936 4.6505
R3000 VDD.n942 VDD.n941 4.6505
R3001 VDD.n947 VDD.n946 4.6505
R3002 VDD.n1018 VDD.n1017 4.6505
R3003 VDD.n878 VDD.n162 4.6505
R3004 VDD.n877 VDD.n876 4.6505
R3005 VDD.n864 VDD.n863 4.6505
R3006 VDD.n859 VDD.n858 4.6505
R3007 VDD.n854 VDD.n853 4.6505
R3008 VDD.n849 VDD.n848 4.6505
R3009 VDD.n844 VDD.n843 4.6505
R3010 VDD.n839 VDD.n838 4.6505
R3011 VDD.n831 VDD.n830 4.6505
R3012 VDD.n826 VDD.n825 4.6505
R3013 VDD.n821 VDD.n820 4.6505
R3014 VDD.n816 VDD.n815 4.6505
R3015 VDD.n811 VDD.n810 4.6505
R3016 VDD.n806 VDD.n805 4.6505
R3017 VDD.n801 VDD.n800 4.6505
R3018 VDD.n796 VDD.n795 4.6505
R3019 VDD.n791 VDD.n790 4.6505
R3020 VDD.n786 VDD.n785 4.6505
R3021 VDD.n781 VDD.n780 4.6505
R3022 VDD.n776 VDD.n775 4.6505
R3023 VDD.n771 VDD.n770 4.6505
R3024 VDD.n766 VDD.n765 4.6505
R3025 VDD.n761 VDD.n760 4.6505
R3026 VDD.n756 VDD.n755 4.6505
R3027 VDD.n751 VDD.n750 4.6505
R3028 VDD.n743 VDD.n742 4.6505
R3029 VDD.n738 VDD.n737 4.6505
R3030 VDD.n733 VDD.n732 4.6505
R3031 VDD.n728 VDD.n727 4.6505
R3032 VDD.n723 VDD.n722 4.6505
R3033 VDD.n718 VDD.n717 4.6505
R3034 VDD.n713 VDD.n712 4.6505
R3035 VDD.n708 VDD.n707 4.6505
R3036 VDD.n703 VDD.n702 4.6505
R3037 VDD.n698 VDD.n697 4.6505
R3038 VDD.n693 VDD.n692 4.6505
R3039 VDD.n688 VDD.n687 4.6505
R3040 VDD.n683 VDD.n682 4.6505
R3041 VDD.n678 VDD.n677 4.6505
R3042 VDD.n673 VDD.n672 4.6505
R3043 VDD.n668 VDD.n667 4.6505
R3044 VDD.n663 VDD.n662 4.6505
R3045 VDD.n655 VDD.n654 4.6505
R3046 VDD.n650 VDD.n649 4.6505
R3047 VDD.n645 VDD.n644 4.6505
R3048 VDD.n640 VDD.n639 4.6505
R3049 VDD.n635 VDD.n634 4.6505
R3050 VDD.n630 VDD.n629 4.6505
R3051 VDD.n625 VDD.n624 4.6505
R3052 VDD.n620 VDD.n619 4.6505
R3053 VDD.n615 VDD.n614 4.6505
R3054 VDD.n610 VDD.n609 4.6505
R3055 VDD.n605 VDD.n604 4.6505
R3056 VDD.n600 VDD.n599 4.6505
R3057 VDD.n595 VDD.n594 4.6505
R3058 VDD.n590 VDD.n589 4.6505
R3059 VDD.n585 VDD.n584 4.6505
R3060 VDD.n580 VDD.n579 4.6505
R3061 VDD.n575 VDD.n574 4.6505
R3062 VDD.n567 VDD.n566 4.6505
R3063 VDD.n562 VDD.n561 4.6505
R3064 VDD.n557 VDD.n556 4.6505
R3065 VDD.n552 VDD.n551 4.6505
R3066 VDD.n547 VDD.n546 4.6505
R3067 VDD.n542 VDD.n541 4.6505
R3068 VDD.n537 VDD.n536 4.6505
R3069 VDD.n532 VDD.n531 4.6505
R3070 VDD.n527 VDD.n526 4.6505
R3071 VDD.n522 VDD.n521 4.6505
R3072 VDD.n517 VDD.n516 4.6505
R3073 VDD.n512 VDD.n511 4.6505
R3074 VDD.n507 VDD.n506 4.6505
R3075 VDD.n502 VDD.n501 4.6505
R3076 VDD.n497 VDD.n496 4.6505
R3077 VDD.n492 VDD.n491 4.6505
R3078 VDD.n487 VDD.n486 4.6505
R3079 VDD.n479 VDD.n478 4.6505
R3080 VDD.n474 VDD.n473 4.6505
R3081 VDD.n469 VDD.n468 4.6505
R3082 VDD.n464 VDD.n463 4.6505
R3083 VDD.n459 VDD.n458 4.6505
R3084 VDD.n454 VDD.n453 4.6505
R3085 VDD.n449 VDD.n448 4.6505
R3086 VDD.n444 VDD.n443 4.6505
R3087 VDD.n439 VDD.n438 4.6505
R3088 VDD.n434 VDD.n433 4.6505
R3089 VDD.n429 VDD.n428 4.6505
R3090 VDD.n424 VDD.n423 4.6505
R3091 VDD.n419 VDD.n418 4.6505
R3092 VDD.n414 VDD.n413 4.6505
R3093 VDD.n409 VDD.n408 4.6505
R3094 VDD.n404 VDD.n403 4.6505
R3095 VDD.n399 VDD.n398 4.6505
R3096 VDD.n391 VDD.n390 4.6505
R3097 VDD.n386 VDD.n385 4.6505
R3098 VDD.n381 VDD.n380 4.6505
R3099 VDD.n376 VDD.n375 4.6505
R3100 VDD.n181 VDD.n180 4.6505
R3101 VDD.n186 VDD.n185 4.6505
R3102 VDD.n191 VDD.n190 4.6505
R3103 VDD.n196 VDD.n195 4.6505
R3104 VDD.n204 VDD.n203 4.6505
R3105 VDD.n209 VDD.n208 4.6505
R3106 VDD.n214 VDD.n213 4.6505
R3107 VDD.n219 VDD.n218 4.6505
R3108 VDD.n224 VDD.n223 4.6505
R3109 VDD.n229 VDD.n228 4.6505
R3110 VDD.n234 VDD.n233 4.6505
R3111 VDD.n239 VDD.n238 4.6505
R3112 VDD.n249 VDD.n248 4.6505
R3113 VDD.n254 VDD.n253 4.6505
R3114 VDD.n259 VDD.n258 4.6505
R3115 VDD.n244 VDD.n243 4.6505
R3116 VDD.n297 VDD.n296 4.6505
R3117 VDD.n302 VDD.n301 4.6505
R3118 VDD.n307 VDD.n306 4.6505
R3119 VDD.n312 VDD.n311 4.6505
R3120 VDD.n317 VDD.n316 4.6505
R3121 VDD.n322 VDD.n321 4.6505
R3122 VDD.n327 VDD.n326 4.6505
R3123 VDD.n332 VDD.n331 4.6505
R3124 VDD.n337 VDD.n336 4.6505
R3125 VDD.n345 VDD.n344 4.6505
R3126 VDD.n350 VDD.n349 4.6505
R3127 VDD.n355 VDD.n354 4.6505
R3128 VDD.n361 VDD.n360 4.6505
R3129 VDD.n367 VDD.n366 4.6505
R3130 VDD.n6431 VDD.n6430 4.6505
R3131 VDD.n6427 VDD.n6426 4.6505
R3132 VDD.n6421 VDD.n6420 4.6505
R3133 VDD.n6415 VDD.n6414 4.6505
R3134 VDD.n6409 VDD.n6408 4.6505
R3135 VDD.n6403 VDD.n6402 4.6505
R3136 VDD.n6397 VDD.n6396 4.6505
R3137 VDD.n6391 VDD.n6390 4.6505
R3138 VDD.n6385 VDD.n6384 4.6505
R3139 VDD.n6379 VDD.n6378 4.6505
R3140 VDD.n6371 VDD.n6370 4.6505
R3141 VDD.n6365 VDD.n6364 4.6505
R3142 VDD.n6357 VDD.n6356 4.6505
R3143 VDD.n6351 VDD.n6350 4.6505
R3144 VDD.n6345 VDD.n6344 4.6505
R3145 VDD.n6339 VDD.n6338 4.6505
R3146 VDD.n6333 VDD.n6332 4.6505
R3147 VDD.n6327 VDD.n6326 4.6505
R3148 VDD.n6321 VDD.n6320 4.6505
R3149 VDD.n6315 VDD.n6314 4.6505
R3150 VDD.n6309 VDD.n6308 4.6505
R3151 VDD.n6303 VDD.n6302 4.6505
R3152 VDD.n6297 VDD.n6296 4.6505
R3153 VDD.n6291 VDD.n6290 4.6505
R3154 VDD.n6285 VDD.n6284 4.6505
R3155 VDD.n6279 VDD.n6278 4.6505
R3156 VDD.n6273 VDD.n6272 4.6505
R3157 VDD.n6505 VDD.n6504 4.6505
R3158 VDD.n6265 VDD.n6264 4.6505
R3159 VDD.n5492 VDD.n5491 4.51815
R3160 VDD.n5485 VDD.n5484 4.51815
R3161 VDD.n5478 VDD.n5477 4.51815
R3162 VDD.n5471 VDD.n5470 4.51815
R3163 VDD.n5464 VDD.n5463 4.51815
R3164 VDD.n5457 VDD.n5456 4.51815
R3165 VDD.n5450 VDD.n5449 4.51815
R3166 VDD.n5443 VDD.n5442 4.51815
R3167 VDD.n5436 VDD.n5435 4.51815
R3168 VDD.n5429 VDD.n5428 4.51815
R3169 VDD.n5422 VDD.n5421 4.51815
R3170 VDD.n5415 VDD.n5414 4.51815
R3171 VDD.n5408 VDD.n5407 4.51815
R3172 VDD.n5401 VDD.n5400 4.51815
R3173 VDD.n5394 VDD.n5393 4.51815
R3174 VDD.n5387 VDD.n5386 4.51815
R3175 VDD.n5380 VDD.n5379 4.51815
R3176 VDD.n5373 VDD.n5372 4.51815
R3177 VDD.n5366 VDD.n5365 4.51815
R3178 VDD.n5359 VDD.n5358 4.51815
R3179 VDD.n5085 VDD.n5084 4.5005
R3180 VDD.n5066 VDD.n5065 4.5005
R3181 VDD.n5046 VDD.n5045 4.5005
R3182 VDD.n5027 VDD.n5026 4.5005
R3183 VDD.n5006 VDD.n5005 4.5005
R3184 VDD.n4984 VDD.n4983 4.5005
R3185 VDD.n4990 VDD.n4989 4.5005
R3186 VDD.n4961 VDD.n4960 4.5005
R3187 VDD.n4966 VDD.n4965 4.5005
R3188 VDD.n4943 VDD.n4942 4.5005
R3189 VDD.n4918 VDD.n4917 4.5005
R3190 VDD.n4901 VDD.n4900 4.5005
R3191 VDD.n4877 VDD.n4876 4.5005
R3192 VDD.n4858 VDD.n4857 4.5005
R3193 VDD.n4817 VDD.n4816 4.5005
R3194 VDD.n4836 VDD.n4835 4.5005
R3195 VDD.n4794 VDD.n4793 4.5005
R3196 VDD.n4810 VDD.n4809 4.5005
R3197 VDD.n4787 VDD.n4786 4.5005
R3198 VDD.n4751 VDD.n4750 4.5005
R3199 VDD.n4732 VDD.n4731 4.5005
R3200 VDD.n4712 VDD.n4711 4.5005
R3201 VDD.n4693 VDD.n4692 4.5005
R3202 VDD.n4673 VDD.n4672 4.5005
R3203 VDD.n4650 VDD.n4649 4.5005
R3204 VDD.n4656 VDD.n4655 4.5005
R3205 VDD.n4627 VDD.n4626 4.5005
R3206 VDD.n4632 VDD.n4631 4.5005
R3207 VDD.n4609 VDD.n4608 4.5005
R3208 VDD.n4589 VDD.n4588 4.5005
R3209 VDD.n4565 VDD.n4564 4.5005
R3210 VDD.n4547 VDD.n4546 4.5005
R3211 VDD.n4508 VDD.n4507 4.5005
R3212 VDD.n4485 VDD.n4484 4.5005
R3213 VDD.n4502 VDD.n4501 4.5005
R3214 VDD.n4462 VDD.n4461 4.5005
R3215 VDD.n4478 VDD.n4477 4.5005
R3216 VDD.n4438 VDD.n4437 4.5005
R3217 VDD.n4421 VDD.n4420 4.5005
R3218 VDD.n4401 VDD.n4400 4.5005
R3219 VDD.n4384 VDD.n4383 4.5005
R3220 VDD.n4368 VDD.n4367 4.5005
R3221 VDD.n4349 VDD.n4348 4.5005
R3222 VDD.n4328 VDD.n4327 4.5005
R3223 VDD.n4334 VDD.n4333 4.5005
R3224 VDD.n4307 VDD.n4306 4.5005
R3225 VDD.n4312 VDD.n4311 4.5005
R3226 VDD.n4294 VDD.n4293 4.5005
R3227 VDD.n4283 VDD.n4282 4.5005
R3228 VDD.n4267 VDD.n4266 4.5005
R3229 VDD.n4236 VDD.n4235 4.5005
R3230 VDD.n4221 VDD.n4220 4.5005
R3231 VDD.n4201 VDD.n4200 4.5005
R3232 VDD.n4180 VDD.n4179 4.5005
R3233 VDD.n4195 VDD.n4194 4.5005
R3234 VDD.n4160 VDD.n4159 4.5005
R3235 VDD.n4154 VDD.n4153 4.5005
R3236 VDD.n4136 VDD.n4135 4.5005
R3237 VDD.n4118 VDD.n4117 4.5005
R3238 VDD.n4099 VDD.n4098 4.5005
R3239 VDD.n4080 VDD.n4079 4.5005
R3240 VDD.n4065 VDD.n4064 4.5005
R3241 VDD.n4046 VDD.n4045 4.5005
R3242 VDD.n4024 VDD.n4023 4.5005
R3243 VDD.n4030 VDD.n4029 4.5005
R3244 VDD.n4001 VDD.n4000 4.5005
R3245 VDD.n4007 VDD.n4006 4.5005
R3246 VDD.n3984 VDD.n3983 4.5005
R3247 VDD.n3973 VDD.n3972 4.5005
R3248 VDD.n3955 VDD.n3954 4.5005
R3249 VDD.n3934 VDD.n3933 4.5005
R3250 VDD.n3900 VDD.n3899 4.5005
R3251 VDD.n3894 VDD.n3893 4.5005
R3252 VDD.n3884 VDD.n3883 4.5005
R3253 VDD.n3855 VDD.n3854 4.5005
R3254 VDD.n3832 VDD.n3831 4.5005
R3255 VDD.n3849 VDD.n3848 4.5005
R3256 VDD.n3826 VDD.n3825 4.5005
R3257 VDD.n3806 VDD.n3805 4.5005
R3258 VDD.n3786 VDD.n3785 4.5005
R3259 VDD.n3766 VDD.n3765 4.5005
R3260 VDD.n3746 VDD.n3745 4.5005
R3261 VDD.n3727 VDD.n3726 4.5005
R3262 VDD.n3707 VDD.n3706 4.5005
R3263 VDD.n3684 VDD.n3683 4.5005
R3264 VDD.n3691 VDD.n3690 4.5005
R3265 VDD.n3661 VDD.n3660 4.5005
R3266 VDD.n3667 VDD.n3666 4.5005
R3267 VDD.n3644 VDD.n3643 4.5005
R3268 VDD.n3634 VDD.n3633 4.5005
R3269 VDD.n3616 VDD.n3615 4.5005
R3270 VDD.n3595 VDD.n3594 4.5005
R3271 VDD.n3575 VDD.n3574 4.5005
R3272 VDD.n3556 VDD.n3555 4.5005
R3273 VDD.n3532 VDD.n3531 4.5005
R3274 VDD.n3518 VDD.n3517 4.5005
R3275 VDD.n3525 VDD.n3524 4.5005
R3276 VDD.n3491 VDD.n3490 4.5005
R3277 VDD.n3512 VDD.n3511 4.5005
R3278 VDD.n3486 VDD.n3485 4.5005
R3279 VDD.n3465 VDD.n3464 4.5005
R3280 VDD.n3445 VDD.n3444 4.5005
R3281 VDD.n3424 VDD.n3423 4.5005
R3282 VDD.n3404 VDD.n3403 4.5005
R3283 VDD.n3019 VDD.n3018 4.5005
R3284 VDD.n3040 VDD.n3039 4.5005
R3285 VDD.n3001 VDD.n3000 4.5005
R3286 VDD.n3046 VDD.n3045 4.5005
R3287 VDD.n5101 VDD.n5100 4.5005
R3288 VDD.n5120 VDD.n5119 4.5005
R3289 VDD.n5127 VDD.n5126 4.5005
R3290 VDD.n5141 VDD.n5140 4.5005
R3291 VDD.n5152 VDD.n5151 4.5005
R3292 VDD.n5269 VDD.n5268 4.5005
R3293 VDD.n105 VDD.n104 4.5005
R3294 VDD.n95 VDD.n94 4.5005
R3295 VDD.n3733 VDD.n3732 4.4805
R3296 VDD.n3745 VDD.n3744 4.4805
R3297 VDD.n4064 VDD.n4063 4.4805
R3298 VDD.n4088 VDD.n4087 4.4805
R3299 VDD.n4098 VDD.n4097 4.4805
R3300 VDD.n4282 VDD.n4281 4.4805
R3301 VDD.n4366 VDD.n4365 4.4805
R3302 VDD.n4410 VDD.n4409 4.4805
R3303 VDD.n4420 VDD.n4419 4.4805
R3304 VDD.n4711 VDD.n4698 4.4805
R3305 VDD.n4700 VDD.n4699 4.4805
R3306 VDD.n4758 VDD.n4757 4.4805
R3307 VDD.n5026 VDD.n5013 4.4805
R3308 VDD.n5065 VDD.n5052 4.4805
R3309 VDD.n5054 VDD.n5053 4.4805
R3310 VDD.n5197 VDD.n5196 4.22272
R3311 VDD.n1191 VDD.n1189 4.20563
R3312 VDD.n169 VDD.n166 4.18959
R3313 VDD.n3483 VDD.n3473 4.1605
R3314 VDD.n3574 VDD.n3573 4.1605
R3315 VDD.n3573 VDD.n3563 4.1605
R3316 VDD.n3847 VDD.n3837 4.1605
R3317 VDD.n3933 VDD.n3932 4.1605
R3318 VDD.n3932 VDD.n3922 4.1605
R3319 VDD.n4135 VDD.n4134 4.1605
R3320 VDD.n4266 VDD.n4265 4.1605
R3321 VDD.n4265 VDD.n4257 4.1605
R3322 VDD.n4524 VDD.n4512 4.1605
R3323 VDD.n4874 VDD.n4864 4.1605
R3324 VDD.n4876 VDD.n4874 4.1605
R3325 VDD.n5119 VDD.n5109 4.1605
R3326 VDD.n1158 VDD.n1155 4.09507
R3327 VDD.n2894 VDD.n2892 4.03915
R3328 VDD.n4191 VDD.t33 4.03915
R3329 VDD.n146 VDD.t23 4.02461
R3330 VDD.n366 VDD.n363 3.95686
R3331 VDD.n3498 VDD.n3497 3.93153
R3332 VDD.n3542 VDD.n3541 3.93153
R3333 VDD.n3862 VDD.n3861 3.93153
R3334 VDD.n3905 VDD.n3904 3.93153
R3335 VDD.n4207 VDD.n4206 3.93153
R3336 VDD.n4241 VDD.n4240 3.93153
R3337 VDD.n4534 VDD.n4533 3.93153
R3338 VDD.n4569 VDD.n4568 3.93153
R3339 VDD.n4886 VDD.n4885 3.93153
R3340 VDD.n4925 VDD.n4924 3.93153
R3341 VDD.n264 VDD.n261 3.87929
R3342 VDD.n4575 VDD.t21 3.85557
R3343 VDD.n3391 VDD.n3390 3.8405
R3344 VDD.n3403 VDD.n3402 3.8405
R3345 VDD.n3726 VDD.n3725 3.8405
R3346 VDD.n3753 VDD.n3752 3.8405
R3347 VDD.n3765 VDD.n3764 3.8405
R3348 VDD.n3972 VDD.n3971 3.8405
R3349 VDD.n4045 VDD.n4044 3.8405
R3350 VDD.n4107 VDD.n4106 3.8405
R3351 VDD.n4117 VDD.n4116 3.8405
R3352 VDD.n4174 VDD.n4165 3.8405
R3353 VDD.n4347 VDD.n4346 3.8405
R3354 VDD.n4428 VDD.n4427 3.8405
R3355 VDD.n4603 VDD.n4602 3.8405
R3356 VDD.n4681 VDD.n4680 3.8405
R3357 VDD.n4775 VDD.n4774 3.8405
R3358 VDD.n5045 VDD.n5032 3.8405
R3359 VDD.n5034 VDD.n5033 3.8405
R3360 VDD.n162 VDD.n161 3.8405
R3361 VDD.n6208 VDD.n6207 3.76521
R3362 VDD.n6201 VDD.n6200 3.76521
R3363 VDD.n6194 VDD.n6193 3.76521
R3364 VDD.n6187 VDD.n6186 3.76521
R3365 VDD.n6180 VDD.n6179 3.76521
R3366 VDD.n6173 VDD.n6172 3.76521
R3367 VDD.n6166 VDD.n6165 3.76521
R3368 VDD.n6159 VDD.n6158 3.76521
R3369 VDD.n6152 VDD.n6151 3.76521
R3370 VDD.n6145 VDD.n6144 3.76521
R3371 VDD.n6138 VDD.n6137 3.76521
R3372 VDD.n6131 VDD.n6130 3.76521
R3373 VDD.n6124 VDD.n6123 3.76521
R3374 VDD.n6117 VDD.n6116 3.76521
R3375 VDD.n6110 VDD.n6109 3.76521
R3376 VDD.n6103 VDD.n6102 3.76521
R3377 VDD.n6096 VDD.n6095 3.76521
R3378 VDD.n6089 VDD.n6088 3.76521
R3379 VDD.n6082 VDD.n6081 3.76521
R3380 VDD.n6075 VDD.n6074 3.76521
R3381 VDD.n5261 VDD.n5200 3.672
R3382 VDD.n896 VDD.n895 3.53932
R3383 VDD.n2998 VDD.n2997 3.52641
R3384 VDD.n3462 VDD.n3452 3.5205
R3385 VDD.n3485 VDD.n3484 3.5205
R3386 VDD.n3555 VDD.n3554 3.5205
R3387 VDD.n3594 VDD.n3593 3.5205
R3388 VDD.n3593 VDD.n3583 3.5205
R3389 VDD.n3805 VDD.n3804 3.5205
R3390 VDD.n3824 VDD.n3814 3.5205
R3391 VDD.n3954 VDD.n3953 3.5205
R3392 VDD.n3953 VDD.n3943 3.5205
R3393 VDD.n4174 VDD.n4164 3.5205
R3394 VDD.n4194 VDD.n4184 3.5205
R3395 VDD.n5140 VDD.n5130 3.5205
R3396 VDD.n5145 VDD.n5144 3.5205
R3397 VDD.n886 VDD.n885 3.46403
R3398 VDD.n6752 VDD.n6749 3.39063
R3399 VDD.n3507 VDD.n3505 3.30485
R3400 VDD.n3546 VDD.n3544 3.30485
R3401 VDD.n3873 VDD.n3871 3.30485
R3402 VDD.n4211 VDD.n4210 3.30485
R3403 VDD.n4541 VDD.n4539 3.30485
R3404 VDD.n4573 VDD.n4571 3.30485
R3405 VDD.n4895 VDD.n4893 3.30485
R3406 VDD.n4929 VDD.n4927 3.30485
R3407 VDD.n5115 VDD.t24 3.30485
R3408 VDD.n1515 VDD.n1428 3.23078
R3409 VDD.n3018 VDD.n3017 3.2005
R3410 VDD.n3411 VDD.n3410 3.2005
R3411 VDD.n3423 VDD.n3422 3.2005
R3412 VDD.n3517 VDD.n3516 3.2005
R3413 VDD.n3633 VDD.n3632 3.2005
R3414 VDD.n3637 VDD.n3636 3.2005
R3415 VDD.n3706 VDD.n3705 3.2005
R3416 VDD.n3773 VDD.n3772 3.2005
R3417 VDD.n3785 VDD.n3784 3.2005
R3418 VDD.n4023 VDD.n4022 3.2005
R3419 VDD.n4125 VDD.n4124 3.2005
R3420 VDD.n4326 VDD.n4325 3.2005
R3421 VDD.n4446 VDD.n4445 3.2005
R3422 VDD.n4671 VDD.n4670 3.2005
R3423 VDD.n4798 VDD.n4797 3.2005
R3424 VDD.n4960 VDD.n4959 3.2005
R3425 VDD.n4980 VDD.n4970 3.2005
R3426 VDD.n4983 VDD.n4982 3.2005
R3427 VDD.n5015 VDD.n5014 3.2005
R3428 VDD.n1372 VDD.n1371 3.2005
R3429 VDD.n2694 VDD.n2693 3.12939
R3430 VDD.n2995 VDD.n2991 3.12127
R3431 VDD.n3871 VDD.t19 3.12127
R3432 VDD.n4059 VDD.n4056 3.12127
R3433 VDD.n4319 VDD.t129 3.12127
R3434 VDD.n4380 VDD.n4377 3.12127
R3435 VDD.n4728 VDD.n4724 3.12127
R3436 VDD.n4975 VDD.t76 3.12127
R3437 VDD.t120 VDD.n5078 3.12127
R3438 VDD.n4912 VDD.n4911 3.03311
R3439 VDD.n4840 VDD.n4839 3.03311
R3440 VDD.n4557 VDD.n4556 3.03311
R3441 VDD.n4528 VDD.n4527 3.03311
R3442 VDD.n4229 VDD.n4228 3.03311
R3443 VDD.n5146 VDD.n5145 3.03311
R3444 VDD.n3877 VDD.n3876 3.03311
R3445 VDD.n4175 VDD.n4174 3.03311
R3446 VDD.n4456 VDD.n4455 3.03311
R3447 VDD.n4769 VDD.n4768 3.03311
R3448 VDD.n6076 VDD.n6075 3.02889
R3449 VDD.n6083 VDD.n6082 3.02889
R3450 VDD.n6090 VDD.n6089 3.02889
R3451 VDD.n6097 VDD.n6096 3.02889
R3452 VDD.n6104 VDD.n6103 3.02889
R3453 VDD.n6111 VDD.n6110 3.02889
R3454 VDD.n6118 VDD.n6117 3.02889
R3455 VDD.n6125 VDD.n6124 3.02889
R3456 VDD.n6132 VDD.n6131 3.02889
R3457 VDD.n6139 VDD.n6138 3.02889
R3458 VDD.n6146 VDD.n6145 3.02889
R3459 VDD.n6153 VDD.n6152 3.02889
R3460 VDD.n6160 VDD.n6159 3.02889
R3461 VDD.n6167 VDD.n6166 3.02889
R3462 VDD.n6174 VDD.n6173 3.02889
R3463 VDD.n6181 VDD.n6180 3.02889
R3464 VDD.n6188 VDD.n6187 3.02889
R3465 VDD.n6195 VDD.n6194 3.02889
R3466 VDD.n6202 VDD.n6201 3.02889
R3467 VDD.n6209 VDD.n6208 3.02889
R3468 VDD.n5897 VDD.n5896 3.02889
R3469 VDD.n5904 VDD.n5903 3.02889
R3470 VDD.n5911 VDD.n5910 3.02889
R3471 VDD.n5918 VDD.n5917 3.02889
R3472 VDD.n5925 VDD.n5924 3.02889
R3473 VDD.n5932 VDD.n5931 3.02889
R3474 VDD.n5939 VDD.n5938 3.02889
R3475 VDD.n5946 VDD.n5945 3.02889
R3476 VDD.n5953 VDD.n5952 3.02889
R3477 VDD.n5960 VDD.n5959 3.02889
R3478 VDD.n5967 VDD.n5966 3.02889
R3479 VDD.n5974 VDD.n5973 3.02889
R3480 VDD.n5981 VDD.n5980 3.02889
R3481 VDD.n5988 VDD.n5987 3.02889
R3482 VDD.n5995 VDD.n5994 3.02889
R3483 VDD.n6002 VDD.n6001 3.02889
R3484 VDD.n6009 VDD.n6008 3.02889
R3485 VDD.n6016 VDD.n6015 3.02889
R3486 VDD.n6023 VDD.n6022 3.02889
R3487 VDD.n6030 VDD.n6029 3.02889
R3488 VDD.n5718 VDD.n5717 3.02889
R3489 VDD.n5725 VDD.n5724 3.02889
R3490 VDD.n5732 VDD.n5731 3.02889
R3491 VDD.n5739 VDD.n5738 3.02889
R3492 VDD.n5746 VDD.n5745 3.02889
R3493 VDD.n5753 VDD.n5752 3.02889
R3494 VDD.n5760 VDD.n5759 3.02889
R3495 VDD.n5767 VDD.n5766 3.02889
R3496 VDD.n5774 VDD.n5773 3.02889
R3497 VDD.n5781 VDD.n5780 3.02889
R3498 VDD.n5788 VDD.n5787 3.02889
R3499 VDD.n5795 VDD.n5794 3.02889
R3500 VDD.n5802 VDD.n5801 3.02889
R3501 VDD.n5809 VDD.n5808 3.02889
R3502 VDD.n5816 VDD.n5815 3.02889
R3503 VDD.n5823 VDD.n5822 3.02889
R3504 VDD.n5830 VDD.n5829 3.02889
R3505 VDD.n5837 VDD.n5836 3.02889
R3506 VDD.n5844 VDD.n5843 3.02889
R3507 VDD.n5851 VDD.n5850 3.02889
R3508 VDD.n5539 VDD.n5538 3.02889
R3509 VDD.n5546 VDD.n5545 3.02889
R3510 VDD.n5553 VDD.n5552 3.02889
R3511 VDD.n5560 VDD.n5559 3.02889
R3512 VDD.n5567 VDD.n5566 3.02889
R3513 VDD.n5574 VDD.n5573 3.02889
R3514 VDD.n5581 VDD.n5580 3.02889
R3515 VDD.n5588 VDD.n5587 3.02889
R3516 VDD.n5595 VDD.n5594 3.02889
R3517 VDD.n5602 VDD.n5601 3.02889
R3518 VDD.n5609 VDD.n5608 3.02889
R3519 VDD.n5616 VDD.n5615 3.02889
R3520 VDD.n5623 VDD.n5622 3.02889
R3521 VDD.n5630 VDD.n5629 3.02889
R3522 VDD.n5637 VDD.n5636 3.02889
R3523 VDD.n5644 VDD.n5643 3.02889
R3524 VDD.n5651 VDD.n5650 3.02889
R3525 VDD.n5658 VDD.n5657 3.02889
R3526 VDD.n5665 VDD.n5664 3.02889
R3527 VDD.n5672 VDD.n5671 3.02889
R3528 VDD.n5360 VDD.n5359 3.02889
R3529 VDD.n5367 VDD.n5366 3.02889
R3530 VDD.n5374 VDD.n5373 3.02889
R3531 VDD.n5381 VDD.n5380 3.02889
R3532 VDD.n5388 VDD.n5387 3.02889
R3533 VDD.n5395 VDD.n5394 3.02889
R3534 VDD.n5402 VDD.n5401 3.02889
R3535 VDD.n5409 VDD.n5408 3.02889
R3536 VDD.n5416 VDD.n5415 3.02889
R3537 VDD.n5423 VDD.n5422 3.02889
R3538 VDD.n5430 VDD.n5429 3.02889
R3539 VDD.n5437 VDD.n5436 3.02889
R3540 VDD.n5444 VDD.n5443 3.02889
R3541 VDD.n5451 VDD.n5450 3.02889
R3542 VDD.n5458 VDD.n5457 3.02889
R3543 VDD.n5465 VDD.n5464 3.02889
R3544 VDD.n5472 VDD.n5471 3.02889
R3545 VDD.n5479 VDD.n5478 3.02889
R3546 VDD.n5486 VDD.n5485 3.02889
R3547 VDD.n5493 VDD.n5492 3.02889
R3548 VDD.n2517 VDD.n2516 3.02889
R3549 VDD.n2524 VDD.n2523 3.02889
R3550 VDD.n2531 VDD.n2530 3.02889
R3551 VDD.n2538 VDD.n2537 3.02889
R3552 VDD.n2545 VDD.n2544 3.02889
R3553 VDD.n2552 VDD.n2551 3.02889
R3554 VDD.n2559 VDD.n2558 3.02889
R3555 VDD.n2566 VDD.n2565 3.02889
R3556 VDD.n2573 VDD.n2572 3.02889
R3557 VDD.n2580 VDD.n2579 3.02889
R3558 VDD.n2587 VDD.n2586 3.02889
R3559 VDD.n2594 VDD.n2593 3.02889
R3560 VDD.n2601 VDD.n2600 3.02889
R3561 VDD.n2608 VDD.n2607 3.02889
R3562 VDD.n2615 VDD.n2614 3.02889
R3563 VDD.n2622 VDD.n2621 3.02889
R3564 VDD.n2629 VDD.n2628 3.02889
R3565 VDD.n2636 VDD.n2635 3.02889
R3566 VDD.n2643 VDD.n2642 3.02889
R3567 VDD.n2650 VDD.n2649 3.02889
R3568 VDD.n2338 VDD.n2337 3.02889
R3569 VDD.n2345 VDD.n2344 3.02889
R3570 VDD.n2352 VDD.n2351 3.02889
R3571 VDD.n2359 VDD.n2358 3.02889
R3572 VDD.n2366 VDD.n2365 3.02889
R3573 VDD.n2373 VDD.n2372 3.02889
R3574 VDD.n2380 VDD.n2379 3.02889
R3575 VDD.n2387 VDD.n2386 3.02889
R3576 VDD.n2394 VDD.n2393 3.02889
R3577 VDD.n2401 VDD.n2400 3.02889
R3578 VDD.n2408 VDD.n2407 3.02889
R3579 VDD.n2415 VDD.n2414 3.02889
R3580 VDD.n2422 VDD.n2421 3.02889
R3581 VDD.n2429 VDD.n2428 3.02889
R3582 VDD.n2436 VDD.n2435 3.02889
R3583 VDD.n2443 VDD.n2442 3.02889
R3584 VDD.n2450 VDD.n2449 3.02889
R3585 VDD.n2457 VDD.n2456 3.02889
R3586 VDD.n2464 VDD.n2463 3.02889
R3587 VDD.n2471 VDD.n2470 3.02889
R3588 VDD.n2159 VDD.n2158 3.02889
R3589 VDD.n2166 VDD.n2165 3.02889
R3590 VDD.n2173 VDD.n2172 3.02889
R3591 VDD.n2180 VDD.n2179 3.02889
R3592 VDD.n2187 VDD.n2186 3.02889
R3593 VDD.n2194 VDD.n2193 3.02889
R3594 VDD.n2201 VDD.n2200 3.02889
R3595 VDD.n2208 VDD.n2207 3.02889
R3596 VDD.n2215 VDD.n2214 3.02889
R3597 VDD.n2222 VDD.n2221 3.02889
R3598 VDD.n2229 VDD.n2228 3.02889
R3599 VDD.n2236 VDD.n2235 3.02889
R3600 VDD.n2243 VDD.n2242 3.02889
R3601 VDD.n2250 VDD.n2249 3.02889
R3602 VDD.n2257 VDD.n2256 3.02889
R3603 VDD.n2264 VDD.n2263 3.02889
R3604 VDD.n2271 VDD.n2270 3.02889
R3605 VDD.n2278 VDD.n2277 3.02889
R3606 VDD.n2285 VDD.n2284 3.02889
R3607 VDD.n2292 VDD.n2291 3.02889
R3608 VDD.n1978 VDD.n1977 3.02889
R3609 VDD.n1985 VDD.n1984 3.02889
R3610 VDD.n1992 VDD.n1991 3.02889
R3611 VDD.n1999 VDD.n1998 3.02889
R3612 VDD.n2006 VDD.n2005 3.02889
R3613 VDD.n2013 VDD.n2012 3.02889
R3614 VDD.n2020 VDD.n2019 3.02889
R3615 VDD.n2027 VDD.n2026 3.02889
R3616 VDD.n2034 VDD.n2033 3.02889
R3617 VDD.n2041 VDD.n2040 3.02889
R3618 VDD.n2048 VDD.n2047 3.02889
R3619 VDD.n2055 VDD.n2054 3.02889
R3620 VDD.n2062 VDD.n2061 3.02889
R3621 VDD.n2069 VDD.n2068 3.02889
R3622 VDD.n2076 VDD.n2075 3.02889
R3623 VDD.n2083 VDD.n2082 3.02889
R3624 VDD.n2090 VDD.n2089 3.02889
R3625 VDD.n2097 VDD.n2096 3.02889
R3626 VDD.n2104 VDD.n2103 3.02889
R3627 VDD.n2111 VDD.n2110 3.02889
R3628 VDD.n1799 VDD.n1798 3.02889
R3629 VDD.n1806 VDD.n1805 3.02889
R3630 VDD.n1813 VDD.n1812 3.02889
R3631 VDD.n1820 VDD.n1819 3.02889
R3632 VDD.n1827 VDD.n1826 3.02889
R3633 VDD.n1834 VDD.n1833 3.02889
R3634 VDD.n1841 VDD.n1840 3.02889
R3635 VDD.n1848 VDD.n1847 3.02889
R3636 VDD.n1855 VDD.n1854 3.02889
R3637 VDD.n1862 VDD.n1861 3.02889
R3638 VDD.n1869 VDD.n1868 3.02889
R3639 VDD.n1876 VDD.n1875 3.02889
R3640 VDD.n1883 VDD.n1882 3.02889
R3641 VDD.n1890 VDD.n1889 3.02889
R3642 VDD.n1897 VDD.n1896 3.02889
R3643 VDD.n1904 VDD.n1903 3.02889
R3644 VDD.n1911 VDD.n1910 3.02889
R3645 VDD.n1918 VDD.n1917 3.02889
R3646 VDD.n1925 VDD.n1924 3.02889
R3647 VDD.n1932 VDD.n1931 3.02889
R3648 VDD.n6029 VDD.n6028 3.01226
R3649 VDD.n6022 VDD.n6021 3.01226
R3650 VDD.n6015 VDD.n6014 3.01226
R3651 VDD.n6008 VDD.n6007 3.01226
R3652 VDD.n6001 VDD.n6000 3.01226
R3653 VDD.n5994 VDD.n5993 3.01226
R3654 VDD.n5987 VDD.n5986 3.01226
R3655 VDD.n5980 VDD.n5979 3.01226
R3656 VDD.n5973 VDD.n5972 3.01226
R3657 VDD.n5966 VDD.n5965 3.01226
R3658 VDD.n5959 VDD.n5958 3.01226
R3659 VDD.n5952 VDD.n5951 3.01226
R3660 VDD.n5945 VDD.n5944 3.01226
R3661 VDD.n5938 VDD.n5937 3.01226
R3662 VDD.n5931 VDD.n5930 3.01226
R3663 VDD.n5924 VDD.n5923 3.01226
R3664 VDD.n5917 VDD.n5916 3.01226
R3665 VDD.n5910 VDD.n5909 3.01226
R3666 VDD.n5903 VDD.n5902 3.01226
R3667 VDD.n5896 VDD.n5895 3.01226
R3668 VDD.n2994 VDD.n2992 2.9377
R3669 VDD.n3034 VDD.n3032 2.9377
R3670 VDD.n3501 VDD.n3500 2.9377
R3671 VDD.n3700 VDD.n3698 2.9377
R3672 VDD.n3721 VDD.n3719 2.9377
R3673 VDD.n3741 VDD.t80 2.9377
R3674 VDD.n3865 VDD.n3864 2.9377
R3675 VDD.n4058 VDD.n4057 2.9377
R3676 VDD.n4075 VDD.n4074 2.9377
R3677 VDD.n4379 VDD.n4378 2.9377
R3678 VDD.n4396 VDD.n4395 2.9377
R3679 VDD.n4727 VDD.n4725 2.9377
R3680 VDD.n4746 VDD.n4744 2.9377
R3681 VDD.n4889 VDD.n4888 2.9377
R3682 VDD.n5081 VDD.n5079 2.9377
R3683 VDD.n5095 VDD.n5094 2.9377
R3684 VDD.n3039 VDD.n3037 2.8805
R3685 VDD.n3442 VDD.n3432 2.8805
R3686 VDD.n3444 VDD.n3442 2.8805
R3687 VDD.n3464 VDD.n3463 2.8805
R3688 VDD.n3615 VDD.n3614 2.8805
R3689 VDD.n3614 VDD.n3604 2.8805
R3690 VDD.n3803 VDD.n3793 2.8805
R3691 VDD.n4152 VDD.n4144 2.8805
R3692 VDD.n4815 VDD.n4814 2.8805
R3693 VDD.n4845 VDD.n4844 2.8805
R3694 VDD.n5004 VDD.n4994 2.8805
R3695 VDD.n5151 VDD.n5149 2.8805
R3696 VDD.n2787 VDD.n2785 2.87311
R3697 VDD.n2832 VDD.n2830 2.87311
R3698 VDD.n1371 VDD.n1367 2.82647
R3699 VDD.n1367 VDD.n1365 2.82647
R3700 VDD.n1365 VDD.n1362 2.82647
R3701 VDD.n1362 VDD.n1360 2.82647
R3702 VDD.n1360 VDD.n1357 2.82647
R3703 VDD.n838 VDD.n834 2.78311
R3704 VDD.n750 VDD.n746 2.78311
R3705 VDD.n662 VDD.n658 2.78311
R3706 VDD.n574 VDD.n570 2.78311
R3707 VDD.n486 VDD.n482 2.78311
R3708 VDD.n398 VDD.n394 2.78311
R3709 VDD.n1104 VDD.n1103 2.76973
R3710 VDD.n2700 VDD.n2699 2.76367
R3711 VDD.n2699 VDD.n2698 2.76367
R3712 VDD.n2698 VDD.n2697 2.76367
R3713 VDD.n3508 VDD.n3503 2.75412
R3714 VDD.n3588 VDD.t29 2.75412
R3715 VDD.n3678 VDD.n3674 2.75412
R3716 VDD.t143 VDD.n3697 2.75412
R3717 VDD.n3874 VDD.n3867 2.75412
R3718 VDD.n3913 VDD.n3912 2.75412
R3719 VDD.n4040 VDD.n4036 2.75412
R3720 VDD.t33 VDD.n4190 2.75412
R3721 VDD.n4212 VDD.n4209 2.75412
R3722 VDD.n4247 VDD.n4246 2.75412
R3723 VDD.n4579 VDD.n4578 2.75412
R3724 VDD.n4708 VDD.n4704 2.75412
R3725 VDD.n4896 VDD.n4891 2.75412
R3726 VDD.n4935 VDD.n4934 2.75412
R3727 VDD.n5062 VDD.n5058 2.75412
R3728 VDD.n1428 VDD.n1424 2.74624
R3729 VDD.n1424 VDD.n1422 2.74624
R3730 VDD.n1422 VDD.n1419 2.74624
R3731 VDD.n1419 VDD.n1417 2.74624
R3732 VDD.n1417 VDD.n1414 2.74624
R3733 VDD.n344 VDD.n343 2.71565
R3734 VDD.n6782 VDD.n6779 2.71203
R3735 VDD.n6779 VDD.n6776 2.71203
R3736 VDD.n6776 VDD.n6773 2.71203
R3737 VDD.n6773 VDD.n6770 2.71203
R3738 VDD.n6770 VDD.n6767 2.71203
R3739 VDD.n6767 VDD.n6764 2.71203
R3740 VDD.n6764 VDD.n6761 2.71203
R3741 VDD.n6761 VDD.n6758 2.71203
R3742 VDD.n6758 VDD.n6755 2.71203
R3743 VDD.n6755 VDD.n6752 2.71203
R3744 VDD.n1104 VDD.n1080 2.70413
R3745 VDD.n203 VDD.n199 2.63808
R3746 VDD.n203 VDD.n202 2.63808
R3747 VDD.n921 VDD.n917 2.63579
R3748 VDD.n838 VDD.n837 2.6241
R3749 VDD.n750 VDD.n749 2.6241
R3750 VDD.n662 VDD.n661 2.6241
R3751 VDD.n574 VDD.n573 2.6241
R3752 VDD.n486 VDD.n485 2.6241
R3753 VDD.n398 VDD.n397 2.6241
R3754 VDD.n6789 VDD.n6786 2.60371
R3755 VDD.n6495 VDD.n6492 2.59871
R3756 VDD.n6497 VDD.n6495 2.59871
R3757 VDD.n5280 VDD.n5278 2.59871
R3758 VDD.n5352 VDD.n5350 2.59871
R3759 VDD.n71 VDD.n69 2.59871
R3760 VDD.n73 VDD.n71 2.59871
R3761 VDD.n75 VDD.n73 2.59871
R3762 VDD.n78 VDD.n75 2.59871
R3763 VDD.n81 VDD.n78 2.59871
R3764 VDD.n6716 VDD.n6713 2.59871
R3765 VDD.n2703 VDD.n2702 2.5774
R3766 VDD.n2705 VDD.n2704 2.5774
R3767 VDD.n2707 VDD.n2706 2.5774
R3768 VDD.n2709 VDD.n2708 2.5774
R3769 VDD.n2711 VDD.n2710 2.5774
R3770 VDD.n2713 VDD.n2712 2.5774
R3771 VDD.n2715 VDD.n2714 2.5774
R3772 VDD.n2717 VDD.n2716 2.5774
R3773 VDD.n2719 VDD.n2718 2.5774
R3774 VDD.n2721 VDD.n2720 2.5774
R3775 VDD.n2723 VDD.n2722 2.5774
R3776 VDD.n2725 VDD.n2724 2.5774
R3777 VDD.n2727 VDD.n2726 2.5774
R3778 VDD.n2729 VDD.n2728 2.5774
R3779 VDD.n2731 VDD.n2730 2.5774
R3780 VDD.n2734 VDD.n2733 2.5774
R3781 VDD.n2737 VDD.n2736 2.5774
R3782 VDD.n2740 VDD.n2739 2.5774
R3783 VDD.n2743 VDD.n2742 2.5774
R3784 VDD.n2746 VDD.n2745 2.5774
R3785 VDD.n2749 VDD.n2748 2.5774
R3786 VDD.n2752 VDD.n2751 2.5774
R3787 VDD.n2755 VDD.n2754 2.5774
R3788 VDD.n2758 VDD.n2757 2.5774
R3789 VDD.n2761 VDD.n2760 2.5774
R3790 VDD.n2764 VDD.n2763 2.5774
R3791 VDD.n2767 VDD.n2766 2.5774
R3792 VDD.n2770 VDD.n2769 2.5774
R3793 VDD.n2773 VDD.n2772 2.5774
R3794 VDD.n2776 VDD.n2775 2.5774
R3795 VDD.n2779 VDD.n2778 2.5774
R3796 VDD.n2783 VDD.n2781 2.5774
R3797 VDD.n3013 VDD.n3011 2.57055
R3798 VDD.n3478 VDD.n3477 2.57055
R3799 VDD.n3552 VDD.t88 2.57055
R3800 VDD.n3677 VDD.n3675 2.57055
R3801 VDD.n3740 VDD.n3738 2.57055
R3802 VDD.n4039 VDD.n4037 2.57055
R3803 VDD.n4093 VDD.n4092 2.57055
R3804 VDD.n4361 VDD.n4360 2.57055
R3805 VDD.n4415 VDD.n4414 2.57055
R3806 VDD.n4517 VDD.n4516 2.57055
R3807 VDD.n4707 VDD.n4705 2.57055
R3808 VDD.n4765 VDD.n4763 2.57055
R3809 VDD.n4853 VDD.t187 2.57055
R3810 VDD.n4869 VDD.n4868 2.57055
R3811 VDD.n5061 VDD.n5059 2.57055
R3812 VDD.n5114 VDD.n5113 2.57055
R3813 VDD.n3045 VDD.n3044 2.5605
R3814 VDD.n3039 VDD.n3038 2.5605
R3815 VDD.n3432 VDD.n3431 2.5605
R3816 VDD.n3444 VDD.n3443 2.5605
R3817 VDD.n3464 VDD.n3462 2.5605
R3818 VDD.n3524 VDD.n3523 2.5605
R3819 VDD.n3531 VDD.n3528 2.5605
R3820 VDD.n3615 VDD.n3602 2.5605
R3821 VDD.n3604 VDD.n3603 2.5605
R3822 VDD.n3683 VDD.n3682 2.5605
R3823 VDD.n3690 VDD.n3689 2.5605
R3824 VDD.n3793 VDD.n3792 2.5605
R3825 VDD.n3854 VDD.n3853 2.5605
R3826 VDD.n3876 VDD.n3860 2.5605
R3827 VDD.n3976 VDD.n3975 2.5605
R3828 VDD.n4000 VDD.n3999 2.5605
R3829 VDD.n4144 VDD.n4143 2.5605
R3830 VDD.n4287 VDD.n4286 2.5605
R3831 VDD.n4305 VDD.n4304 2.5605
R3832 VDD.n4466 VDD.n4465 2.5605
R3833 VDD.n4646 VDD.n4636 2.5605
R3834 VDD.n4648 VDD.n4647 2.5605
R3835 VDD.n4821 VDD.n4820 2.5605
R3836 VDD.n4994 VDD.n4993 2.5605
R3837 VDD.n344 VDD.n340 2.5605
R3838 VDD.n921 VDD.n920 2.48521
R3839 VDD.n843 VDD.n842 2.4651
R3840 VDD.n755 VDD.n754 2.4651
R3841 VDD.n667 VDD.n666 2.4651
R3842 VDD.n579 VDD.n578 2.4651
R3843 VDD.n491 VDD.n490 2.4651
R3844 VDD.n403 VDD.n402 2.4651
R3845 VDD.n1188 VDD.n1185 2.4386
R3846 VDD.n1185 VDD.n1182 2.4386
R3847 VDD.n1182 VDD.n1179 2.4386
R3848 VDD.n1179 VDD.n1176 2.4386
R3849 VDD.n1176 VDD.n1173 2.4386
R3850 VDD.n1173 VDD.n1170 2.4386
R3851 VDD.n1170 VDD.n1167 2.4386
R3852 VDD.n1167 VDD.n1164 2.4386
R3853 VDD.n1164 VDD.n1161 2.4386
R3854 VDD.n1161 VDD.n1158 2.4386
R3855 VDD.n6501 VDD.n6498 2.40766
R3856 VDD.n349 VDD.n348 2.40535
R3857 VDD.n3481 VDD.n3480 2.38697
R3858 VDD.n3571 VDD.n3570 2.38697
R3859 VDD.n3654 VDD.n3650 2.38697
R3860 VDD.t0 VDD.n3841 2.38697
R3861 VDD.n3845 VDD.n3844 2.38697
R3862 VDD.n3930 VDD.n3929 2.38697
R3863 VDD.n4018 VDD.n4014 2.38697
R3864 VDD.n4073 VDD.t47 2.38697
R3865 VDD.n4191 VDD.n4189 2.38697
R3866 VDD.n4263 VDD.n4262 2.38697
R3867 VDD.n4343 VDD.n4340 2.38697
R3868 VDD.n4522 VDD.n4519 2.38697
R3869 VDD.n4597 VDD.n4596 2.38697
R3870 VDD.n4689 VDD.n4685 2.38697
R3871 VDD.n4705 VDD.t15 2.38697
R3872 VDD.n4872 VDD.n4871 2.38697
R3873 VDD.n4955 VDD.n4954 2.38697
R3874 VDD.n5042 VDD.n5038 2.38697
R3875 VDD.n2701 VDD.n2694 2.35733
R3876 VDD.n926 VDD.n925 2.33462
R3877 VDD.n5276 VDD.n5274 2.33125
R3878 VDD.n195 VDD.n194 2.32777
R3879 VDD.n208 VDD.n207 2.32777
R3880 VDD.n830 VDD.n829 2.30609
R3881 VDD.n742 VDD.n741 2.30609
R3882 VDD.n654 VDD.n653 2.30609
R3883 VDD.n566 VDD.n565 2.30609
R3884 VDD.n478 VDD.n477 2.30609
R3885 VDD.n390 VDD.n389 2.30609
R3886 VDD.n5850 VDD.n5849 2.25932
R3887 VDD.n5843 VDD.n5842 2.25932
R3888 VDD.n5836 VDD.n5835 2.25932
R3889 VDD.n5829 VDD.n5828 2.25932
R3890 VDD.n5822 VDD.n5821 2.25932
R3891 VDD.n5815 VDD.n5814 2.25932
R3892 VDD.n5808 VDD.n5807 2.25932
R3893 VDD.n5801 VDD.n5800 2.25932
R3894 VDD.n5794 VDD.n5793 2.25932
R3895 VDD.n5787 VDD.n5786 2.25932
R3896 VDD.n5780 VDD.n5779 2.25932
R3897 VDD.n5773 VDD.n5772 2.25932
R3898 VDD.n5766 VDD.n5765 2.25932
R3899 VDD.n5759 VDD.n5758 2.25932
R3900 VDD.n5752 VDD.n5751 2.25932
R3901 VDD.n5745 VDD.n5744 2.25932
R3902 VDD.n5738 VDD.n5737 2.25932
R3903 VDD.n5731 VDD.n5730 2.25932
R3904 VDD.n5724 VDD.n5723 2.25932
R3905 VDD.n5717 VDD.n5716 2.25932
R3906 VDD.n5671 VDD.n5670 2.25932
R3907 VDD.n5664 VDD.n5663 2.25932
R3908 VDD.n5657 VDD.n5656 2.25932
R3909 VDD.n5650 VDD.n5649 2.25932
R3910 VDD.n5643 VDD.n5642 2.25932
R3911 VDD.n5636 VDD.n5635 2.25932
R3912 VDD.n5629 VDD.n5628 2.25932
R3913 VDD.n5622 VDD.n5621 2.25932
R3914 VDD.n5615 VDD.n5614 2.25932
R3915 VDD.n5608 VDD.n5607 2.25932
R3916 VDD.n5601 VDD.n5600 2.25932
R3917 VDD.n5594 VDD.n5593 2.25932
R3918 VDD.n5587 VDD.n5586 2.25932
R3919 VDD.n5580 VDD.n5579 2.25932
R3920 VDD.n5573 VDD.n5572 2.25932
R3921 VDD.n5566 VDD.n5565 2.25932
R3922 VDD.n5559 VDD.n5558 2.25932
R3923 VDD.n5552 VDD.n5551 2.25932
R3924 VDD.n5545 VDD.n5544 2.25932
R3925 VDD.n5538 VDD.n5537 2.25932
R3926 VDD.n1931 VDD.n1930 2.25932
R3927 VDD.n1924 VDD.n1923 2.25932
R3928 VDD.n1917 VDD.n1916 2.25932
R3929 VDD.n1910 VDD.n1909 2.25932
R3930 VDD.n1903 VDD.n1902 2.25932
R3931 VDD.n1896 VDD.n1895 2.25932
R3932 VDD.n1889 VDD.n1888 2.25932
R3933 VDD.n1882 VDD.n1881 2.25932
R3934 VDD.n1875 VDD.n1874 2.25932
R3935 VDD.n1868 VDD.n1867 2.25932
R3936 VDD.n1861 VDD.n1860 2.25932
R3937 VDD.n1854 VDD.n1853 2.25932
R3938 VDD.n1847 VDD.n1846 2.25932
R3939 VDD.n1840 VDD.n1839 2.25932
R3940 VDD.n1833 VDD.n1832 2.25932
R3941 VDD.n1826 VDD.n1825 2.25932
R3942 VDD.n1819 VDD.n1818 2.25932
R3943 VDD.n1812 VDD.n1811 2.25932
R3944 VDD.n1805 VDD.n1804 2.25932
R3945 VDD.n1798 VDD.n1797 2.25932
R3946 VDD.n131 VDD.n128 2.25932
R3947 VDD.n119 VDD.n116 2.25932
R3948 VDD.n336 VDD.n335 2.2502
R3949 VDD.n3022 VDD.n3021 2.2405
R3950 VDD.n3018 VDD.n3016 2.2405
R3951 VDD.n3421 VDD.n3411 2.2405
R3952 VDD.n3423 VDD.n3421 2.2405
R3953 VDD.n3490 VDD.n3489 2.2405
R3954 VDD.n3633 VDD.n3622 2.2405
R3955 VDD.n3783 VDD.n3773 2.2405
R3956 VDD.n3785 VDD.n3783 2.2405
R3957 VDD.n3831 VDD.n3830 2.2405
R3958 VDD.n4028 VDD.n4027 2.2405
R3959 VDD.n4133 VDD.n4125 2.2405
R3960 VDD.n4159 VDD.n4158 2.2405
R3961 VDD.n4455 VDD.n4446 2.2405
R3962 VDD.n4477 VDD.n4466 2.2405
R3963 VDD.n4483 VDD.n4482 2.2405
R3964 VDD.n4501 VDD.n4489 2.2405
R3965 VDD.n4989 VDD.n4988 2.2405
R3966 VDD.n5025 VDD.n5015 2.2405
R3967 VDD.n2989 VDD.n2987 2.2034
R3968 VDD.n3398 VDD.n3396 2.2034
R3969 VDD.n3457 VDD.n3456 2.2034
R3970 VDD.n3460 VDD.t42 2.2034
R3971 VDD.n3653 VDD.n3651 2.2034
R3972 VDD.n3760 VDD.n3758 2.2034
R3973 VDD.n3819 VDD.n3818 2.2034
R3974 VDD.n4017 VDD.n4015 2.2034
R3975 VDD.n4169 VDD.n4168 2.2034
R3976 VDD.n4342 VDD.n4341 2.2034
R3977 VDD.n4433 VDD.n4432 2.2034
R3978 VDD.n4688 VDD.n4686 2.2034
R3979 VDD.n4782 VDD.n4780 2.2034
R3980 VDD.n5041 VDD.n5039 2.2034
R3981 VDD.n5135 VDD.n5134 2.2034
R3982 VDD.n913 VDD.n912 2.18403
R3983 VDD.n1189 VDD.n1188 2.15176
R3984 VDD.n848 VDD.n847 2.14708
R3985 VDD.n760 VDD.n759 2.14708
R3986 VDD.n672 VDD.n671 2.14708
R3987 VDD.n584 VDD.n583 2.14708
R3988 VDD.n496 VDD.n495 2.14708
R3989 VDD.n408 VDD.n407 2.14708
R3990 VDD.n6504 VDD.n6501 2.10199
R3991 VDD.n354 VDD.n353 2.09505
R3992 VDD.n931 VDD.n930 2.03344
R3993 VDD.n2696 VDD.n2695 2.03225
R3994 VDD.n6507 VDD.n6506 2.03225
R3995 VDD.n6509 VDD.n6508 2.03225
R3996 VDD.n6511 VDD.n6510 2.03225
R3997 VDD.n6513 VDD.n6512 2.03225
R3998 VDD.n6515 VDD.n6514 2.03225
R3999 VDD.n6517 VDD.n6516 2.03225
R4000 VDD.n6519 VDD.n6518 2.03225
R4001 VDD.n6521 VDD.n6520 2.03225
R4002 VDD.n6523 VDD.n6522 2.03225
R4003 VDD.n6525 VDD.n6524 2.03225
R4004 VDD.n6527 VDD.n6526 2.03225
R4005 VDD.n6529 VDD.n6528 2.03225
R4006 VDD.n6531 VDD.n6530 2.03225
R4007 VDD.n6533 VDD.n6532 2.03225
R4008 VDD.n6535 VDD.n6534 2.03225
R4009 VDD.n6537 VDD.n6536 2.03225
R4010 VDD.n6539 VDD.n6538 2.03225
R4011 VDD.n6541 VDD.n6540 2.03225
R4012 VDD.n6543 VDD.n6542 2.03225
R4013 VDD.n6545 VDD.n6544 2.03225
R4014 VDD.n6547 VDD.n6546 2.03225
R4015 VDD.n6549 VDD.n6548 2.03225
R4016 VDD.n6551 VDD.n6550 2.03225
R4017 VDD.n6553 VDD.n6552 2.03225
R4018 VDD.n6555 VDD.n6554 2.03225
R4019 VDD.n6557 VDD.n6556 2.03225
R4020 VDD.n6559 VDD.n6558 2.03225
R4021 VDD.n6561 VDD.n6560 2.03225
R4022 VDD.n6563 VDD.n6562 2.03225
R4023 VDD.n6565 VDD.n6564 2.03225
R4024 VDD.n6567 VDD.n6566 2.03225
R4025 VDD.n6569 VDD.n6568 2.03225
R4026 VDD.n6571 VDD.n6570 2.03225
R4027 VDD.n6574 VDD.n6572 2.03225
R4028 VDD.n6577 VDD.n6575 2.03225
R4029 VDD.n6581 VDD.n6579 2.03225
R4030 VDD.n6585 VDD.n6583 2.03225
R4031 VDD.n6589 VDD.n6587 2.03225
R4032 VDD.n6593 VDD.n6591 2.03225
R4033 VDD.n6597 VDD.n6595 2.03225
R4034 VDD.n6601 VDD.n6599 2.03225
R4035 VDD.n6605 VDD.n6603 2.03225
R4036 VDD.n6609 VDD.n6607 2.03225
R4037 VDD.n6613 VDD.n6611 2.03225
R4038 VDD.n6617 VDD.n6615 2.03225
R4039 VDD.n6621 VDD.n6619 2.03225
R4040 VDD.n6695 VDD.n6693 2.03225
R4041 VDD.n6691 VDD.n6689 2.03225
R4042 VDD.n6687 VDD.n6685 2.03225
R4043 VDD.n6683 VDD.n6681 2.03225
R4044 VDD.n6679 VDD.n6677 2.03225
R4045 VDD.n6675 VDD.n6673 2.03225
R4046 VDD.n6671 VDD.n6669 2.03225
R4047 VDD.n6667 VDD.n6665 2.03225
R4048 VDD.n6663 VDD.n6661 2.03225
R4049 VDD.n6659 VDD.n6657 2.03225
R4050 VDD.n6655 VDD.n6653 2.03225
R4051 VDD.n6651 VDD.n6650 2.03225
R4052 VDD.n6649 VDD.n6648 2.03225
R4053 VDD.n6647 VDD.n6646 2.03225
R4054 VDD.n6645 VDD.n6644 2.03225
R4055 VDD.n6643 VDD.n6642 2.03225
R4056 VDD.n6641 VDD.n6640 2.03225
R4057 VDD.n6639 VDD.n6638 2.03225
R4058 VDD.n6637 VDD.n6636 2.03225
R4059 VDD.n6635 VDD.n6634 2.03225
R4060 VDD.n6633 VDD.n6632 2.03225
R4061 VDD.n6631 VDD.n6630 2.03225
R4062 VDD.n6629 VDD.n6628 2.03225
R4063 VDD.n6627 VDD.n6626 2.03225
R4064 VDD.n6625 VDD.n6624 2.03225
R4065 VDD.n6623 VDD.n6622 2.03225
R4066 VDD.n6433 VDD.n6432 2.03225
R4067 VDD.n6435 VDD.n6434 2.03225
R4068 VDD.n6437 VDD.n6436 2.03225
R4069 VDD.n6439 VDD.n6438 2.03225
R4070 VDD.n6441 VDD.n6440 2.03225
R4071 VDD.n6443 VDD.n6442 2.03225
R4072 VDD.n6445 VDD.n6444 2.03225
R4073 VDD.n6447 VDD.n6446 2.03225
R4074 VDD.n6449 VDD.n6448 2.03225
R4075 VDD.n6451 VDD.n6450 2.03225
R4076 VDD.n6453 VDD.n6452 2.03225
R4077 VDD.n6455 VDD.n6454 2.03225
R4078 VDD.n6457 VDD.n6456 2.03225
R4079 VDD.n6459 VDD.n6458 2.03225
R4080 VDD.n6461 VDD.n6460 2.03225
R4081 VDD.n6463 VDD.n6462 2.03225
R4082 VDD.n6466 VDD.n6464 2.03225
R4083 VDD.n6469 VDD.n6467 2.03225
R4084 VDD.n6473 VDD.n6471 2.03225
R4085 VDD.n6477 VDD.n6475 2.03225
R4086 VDD.n6481 VDD.n6479 2.03225
R4087 VDD.n6485 VDD.n6483 2.03225
R4088 VDD.n3460 VDD.n3459 2.01982
R4089 VDD.n3591 VDD.n3590 2.01982
R4090 VDD.n3630 VDD.n3626 2.01982
R4091 VDD.n3822 VDD.n3821 2.01982
R4092 VDD.n3926 VDD.t91 2.01982
R4093 VDD.n3951 VDD.n3950 2.01982
R4094 VDD.n3994 VDD.n3990 2.01982
R4095 VDD.n4172 VDD.n4170 2.01982
R4096 VDD.n4243 VDD.t105 2.01982
R4097 VDD.n4279 VDD.n4278 2.01982
R4098 VDD.n4322 VDD.n4319 2.01982
R4099 VDD.n4498 VDD.n4497 2.01982
R4100 VDD.n4621 VDD.n4620 2.01982
R4101 VDD.n4667 VDD.n4663 2.01982
R4102 VDD.n4853 VDD.n4852 2.01982
R4103 VDD.n4978 VDD.n4977 2.01982
R4104 VDD.n5023 VDD.n5019 2.01982
R4105 VDD.n190 VDD.n189 2.01747
R4106 VDD.n213 VDD.n212 2.01747
R4107 VDD.n825 VDD.n824 1.98808
R4108 VDD.n737 VDD.n736 1.98808
R4109 VDD.n649 VDD.n648 1.98808
R4110 VDD.n561 VDD.n560 1.98808
R4111 VDD.n473 VDD.n472 1.98808
R4112 VDD.n385 VDD.n384 1.98808
R4113 VDD.n2996 VDD.n2837 1.96602
R4114 VDD.n3036 VDD.n3029 1.96602
R4115 VDD.n3702 VDD.n3695 1.96602
R4116 VDD.n3723 VDD.n3716 1.96602
R4117 VDD.n4060 VDD.n4055 1.96602
R4118 VDD.n4077 VDD.n4072 1.96602
R4119 VDD.n4381 VDD.n4376 1.96602
R4120 VDD.n4398 VDD.n4393 1.96602
R4121 VDD.n4729 VDD.n4722 1.96602
R4122 VDD.n4748 VDD.n4741 1.96602
R4123 VDD.n5082 VDD.n5077 1.96602
R4124 VDD.n5097 VDD.n5092 1.96602
R4125 VDD.n331 VDD.n330 1.93989
R4126 VDD.n3000 VDD.n2999 1.9205
R4127 VDD.n3452 VDD.n3451 1.9205
R4128 VDD.n3485 VDD.n3483 1.9205
R4129 VDD.n3555 VDD.n3538 1.9205
R4130 VDD.n3594 VDD.n3581 1.9205
R4131 VDD.n3583 VDD.n3582 1.9205
R4132 VDD.n3660 VDD.n3658 1.9205
R4133 VDD.n3660 VDD.n3659 1.9205
R4134 VDD.n3683 VDD.n3681 1.9205
R4135 VDD.n3706 VDD.n3704 1.9205
R4136 VDD.n3805 VDD.n3803 1.9205
R4137 VDD.n3814 VDD.n3813 1.9205
R4138 VDD.n3883 VDD.n3880 1.9205
R4139 VDD.n3954 VDD.n3941 1.9205
R4140 VDD.n3943 VDD.n3942 1.9205
R4141 VDD.n4164 VDD.n4163 1.9205
R4142 VDD.n4179 VDD.n4178 1.9205
R4143 VDD.n4193 VDD.n4185 1.9205
R4144 VDD.n4286 VDD.n4285 1.9205
R4145 VDD.n4324 VDD.n4316 1.9205
R4146 VDD.n4461 VDD.n4460 1.9205
R4147 VDD.n4489 VDD.n4488 1.9205
R4148 VDD.n4626 VDD.n4625 1.9205
R4149 VDD.n4625 VDD.n4624 1.9205
R4150 VDD.n4649 VDD.n4648 1.9205
R4151 VDD.n4672 VDD.n4671 1.9205
R4152 VDD.n4835 VDD.n4834 1.9205
R4153 VDD.n4844 VDD.n4843 1.9205
R4154 VDD.n4982 VDD.n4981 1.9205
R4155 VDD.n2833 VDD.n2787 1.90149
R4156 VDD.n2291 VDD.n2290 1.88285
R4157 VDD.n2284 VDD.n2283 1.88285
R4158 VDD.n2277 VDD.n2276 1.88285
R4159 VDD.n2270 VDD.n2269 1.88285
R4160 VDD.n2263 VDD.n2262 1.88285
R4161 VDD.n2256 VDD.n2255 1.88285
R4162 VDD.n2249 VDD.n2248 1.88285
R4163 VDD.n2242 VDD.n2241 1.88285
R4164 VDD.n2235 VDD.n2234 1.88285
R4165 VDD.n2228 VDD.n2227 1.88285
R4166 VDD.n2221 VDD.n2220 1.88285
R4167 VDD.n2214 VDD.n2213 1.88285
R4168 VDD.n2207 VDD.n2206 1.88285
R4169 VDD.n2200 VDD.n2199 1.88285
R4170 VDD.n2193 VDD.n2192 1.88285
R4171 VDD.n2186 VDD.n2185 1.88285
R4172 VDD.n2179 VDD.n2178 1.88285
R4173 VDD.n2172 VDD.n2171 1.88285
R4174 VDD.n2165 VDD.n2164 1.88285
R4175 VDD.n2158 VDD.n2157 1.88285
R4176 VDD.n2110 VDD.n2109 1.88285
R4177 VDD.n2103 VDD.n2102 1.88285
R4178 VDD.n2096 VDD.n2095 1.88285
R4179 VDD.n2089 VDD.n2088 1.88285
R4180 VDD.n2082 VDD.n2081 1.88285
R4181 VDD.n2075 VDD.n2074 1.88285
R4182 VDD.n2068 VDD.n2067 1.88285
R4183 VDD.n2061 VDD.n2060 1.88285
R4184 VDD.n2054 VDD.n2053 1.88285
R4185 VDD.n2047 VDD.n2046 1.88285
R4186 VDD.n2040 VDD.n2039 1.88285
R4187 VDD.n2033 VDD.n2032 1.88285
R4188 VDD.n2026 VDD.n2025 1.88285
R4189 VDD.n2019 VDD.n2018 1.88285
R4190 VDD.n2012 VDD.n2011 1.88285
R4191 VDD.n2005 VDD.n2004 1.88285
R4192 VDD.n1998 VDD.n1997 1.88285
R4193 VDD.n1991 VDD.n1990 1.88285
R4194 VDD.n1984 VDD.n1983 1.88285
R4195 VDD.n1977 VDD.n1976 1.88285
R4196 VDD.n908 VDD.n907 1.88285
R4197 VDD.n3418 VDD.n3416 1.83625
R4198 VDD.n3437 VDD.n3436 1.83625
R4199 VDD.n3629 VDD.n3627 1.83625
R4200 VDD.n3780 VDD.n3778 1.83625
R4201 VDD.n3798 VDD.n3797 1.83625
R4202 VDD.n3993 VDD.n3991 1.83625
R4203 VDD.n4130 VDD.n4129 1.83625
R4204 VDD.n4148 VDD.n4147 1.83625
R4205 VDD.n4321 VDD.n4320 1.83625
R4206 VDD.n4362 VDD.t78 1.83625
R4207 VDD.n4452 VDD.n4450 1.83625
R4208 VDD.n4471 VDD.n4470 1.83625
R4209 VDD.n4805 VDD.n4803 1.83625
R4210 VDD.n4827 VDD.n4826 1.83625
R4211 VDD.n5022 VDD.n5020 1.83625
R4212 VDD.n5158 VDD.n5157 1.83625
R4213 VDD.n853 VDD.n852 1.82907
R4214 VDD.n765 VDD.n764 1.82907
R4215 VDD.n677 VDD.n676 1.82907
R4216 VDD.n589 VDD.n588 1.82907
R4217 VDD.n501 VDD.n500 1.82907
R4218 VDD.n413 VDD.n412 1.82907
R4219 VDD.n360 VDD.n359 1.78474
R4220 VDD.n2702 VDD.n2701 1.77476
R4221 VDD.n936 VDD.n935 1.73226
R4222 VDD.n5353 VDD.n5280 1.7199
R4223 VDD.n185 VDD.n184 1.70717
R4224 VDD.n218 VDD.n217 1.70717
R4225 VDD.n87 VDD.n85 1.69185
R4226 VDD.n6790 VDD.n6716 1.68169
R4227 VDD.n820 VDD.n819 1.67007
R4228 VDD.n732 VDD.n731 1.67007
R4229 VDD.n644 VDD.n643 1.67007
R4230 VDD.n556 VDD.n555 1.67007
R4231 VDD.n468 VDD.n467 1.67007
R4232 VDD.n380 VDD.n379 1.67007
R4233 VDD.n889 VDD.n886 1.65697
R4234 VDD.n3440 VDD.n3439 1.65267
R4235 VDD.n3612 VDD.n3608 1.65267
R4236 VDD.n3612 VDD.n3611 1.65267
R4237 VDD.n3797 VDD.t4 1.65267
R4238 VDD.n3801 VDD.n3800 1.65267
R4239 VDD.n3969 VDD.n3965 1.65267
R4240 VDD.n4112 VDD.t135 1.65267
R4241 VDD.n4150 VDD.n4149 1.65267
R4242 VDD.n4300 VDD.n4297 1.65267
R4243 VDD.n4300 VDD.n4299 1.65267
R4244 VDD.n4474 VDD.n4473 1.65267
R4245 VDD.n4495 VDD.t110 1.65267
R4246 VDD.n4644 VDD.n4640 1.65267
R4247 VDD.n4644 VDD.n4643 1.65267
R4248 VDD.n4832 VDD.n4829 1.65267
R4249 VDD.n5002 VDD.n4998 1.65267
R4250 VDD.n5002 VDD.n5001 1.65267
R4251 VDD.n2828 VDD.n2826 1.64802
R4252 VDD.n2824 VDD.n2823 1.64802
R4253 VDD.n2821 VDD.n2820 1.64802
R4254 VDD.n2818 VDD.n2817 1.64802
R4255 VDD.n2815 VDD.n2814 1.64802
R4256 VDD.n2812 VDD.n2811 1.64802
R4257 VDD.n2809 VDD.n2808 1.64802
R4258 VDD.n2806 VDD.n2805 1.64802
R4259 VDD.n2803 VDD.n2802 1.64802
R4260 VDD.n2800 VDD.n2799 1.64802
R4261 VDD.n2797 VDD.n2796 1.64802
R4262 VDD.n2794 VDD.n2793 1.64802
R4263 VDD.n2791 VDD.n2790 1.64802
R4264 VDD.n1023 VDD.n1021 1.64802
R4265 VDD.n1026 VDD.n1024 1.64802
R4266 VDD.n1029 VDD.n1027 1.64802
R4267 VDD.n1032 VDD.n1030 1.64802
R4268 VDD.n1035 VDD.n1033 1.64802
R4269 VDD.n1038 VDD.n1036 1.64802
R4270 VDD.n1041 VDD.n1039 1.64802
R4271 VDD.n1044 VDD.n1042 1.64802
R4272 VDD.n1047 VDD.n1045 1.64802
R4273 VDD.n1050 VDD.n1048 1.64802
R4274 VDD.n1053 VDD.n1051 1.64802
R4275 VDD.n1056 VDD.n1054 1.64802
R4276 VDD.n1060 VDD.n1058 1.64802
R4277 VDD.n1064 VDD.n1062 1.64802
R4278 VDD.n1068 VDD.n1066 1.64802
R4279 VDD.n1072 VDD.n1070 1.64802
R4280 VDD.n1076 VDD.n1074 1.64802
R4281 VDD.n1080 VDD.n1078 1.64802
R4282 VDD.n326 VDD.n325 1.62959
R4283 VDD.n3401 VDD.n3391 1.6005
R4284 VDD.n3403 VDD.n3401 1.6005
R4285 VDD.n3643 VDD.n3642 1.6005
R4286 VDD.n3711 VDD.n3710 1.6005
R4287 VDD.n3726 VDD.n3724 1.6005
R4288 VDD.n3763 VDD.n3753 1.6005
R4289 VDD.n3765 VDD.n3763 1.6005
R4290 VDD.n3972 VDD.n3961 1.6005
R4291 VDD.n3998 VDD.n3997 1.6005
R4292 VDD.n4021 VDD.n4020 1.6005
R4293 VDD.n4115 VDD.n4107 1.6005
R4294 VDD.n4117 VDD.n4115 1.6005
R4295 VDD.n4327 VDD.n4324 1.6005
R4296 VDD.n4332 VDD.n4331 1.6005
R4297 VDD.n4436 VDD.n4428 1.6005
R4298 VDD.n4626 VDD.n4623 1.6005
R4299 VDD.n4655 VDD.n4654 1.6005
R4300 VDD.n4691 VDD.n4681 1.6005
R4301 VDD.n4965 VDD.n4964 1.6005
R4302 VDD.n5045 VDD.n5044 1.6005
R4303 VDD.n5044 VDD.n5034 1.6005
R4304 VDD.n5125 VDD.n5124 1.6005
R4305 VDD.n5139 VDD.n5138 1.6005
R4306 VDD.n899 VDD.n896 1.58168
R4307 VDD.n858 VDD.n857 1.51106
R4308 VDD.n770 VDD.n769 1.51106
R4309 VDD.n682 VDD.n681 1.51106
R4310 VDD.n594 VDD.n593 1.51106
R4311 VDD.n506 VDD.n505 1.51106
R4312 VDD.n418 VDD.n417 1.51106
R4313 VDD.n2649 VDD.n2648 1.50638
R4314 VDD.n2642 VDD.n2641 1.50638
R4315 VDD.n2635 VDD.n2634 1.50638
R4316 VDD.n2628 VDD.n2627 1.50638
R4317 VDD.n2621 VDD.n2620 1.50638
R4318 VDD.n2614 VDD.n2613 1.50638
R4319 VDD.n2607 VDD.n2606 1.50638
R4320 VDD.n2600 VDD.n2599 1.50638
R4321 VDD.n2593 VDD.n2592 1.50638
R4322 VDD.n2586 VDD.n2585 1.50638
R4323 VDD.n2579 VDD.n2578 1.50638
R4324 VDD.n2572 VDD.n2571 1.50638
R4325 VDD.n2565 VDD.n2564 1.50638
R4326 VDD.n2558 VDD.n2557 1.50638
R4327 VDD.n2551 VDD.n2550 1.50638
R4328 VDD.n2544 VDD.n2543 1.50638
R4329 VDD.n2537 VDD.n2536 1.50638
R4330 VDD.n2530 VDD.n2529 1.50638
R4331 VDD.n2523 VDD.n2522 1.50638
R4332 VDD.n2516 VDD.n2515 1.50638
R4333 VDD.n2470 VDD.n2469 1.50638
R4334 VDD.n2463 VDD.n2462 1.50638
R4335 VDD.n2456 VDD.n2455 1.50638
R4336 VDD.n2449 VDD.n2448 1.50638
R4337 VDD.n2442 VDD.n2441 1.50638
R4338 VDD.n2435 VDD.n2434 1.50638
R4339 VDD.n2428 VDD.n2427 1.50638
R4340 VDD.n2421 VDD.n2420 1.50638
R4341 VDD.n2414 VDD.n2413 1.50638
R4342 VDD.n2407 VDD.n2406 1.50638
R4343 VDD.n2400 VDD.n2399 1.50638
R4344 VDD.n2393 VDD.n2392 1.50638
R4345 VDD.n2386 VDD.n2385 1.50638
R4346 VDD.n2379 VDD.n2378 1.50638
R4347 VDD.n2372 VDD.n2371 1.50638
R4348 VDD.n2365 VDD.n2364 1.50638
R4349 VDD.n2358 VDD.n2357 1.50638
R4350 VDD.n2351 VDD.n2350 1.50638
R4351 VDD.n2344 VDD.n2343 1.50638
R4352 VDD.n2337 VDD.n2336 1.50638
R4353 VDD.n5356 VDD.n5355 1.5005
R4354 VDD.n5348 VDD.n5346 1.49065
R4355 VDD.n5344 VDD.n5342 1.49065
R4356 VDD.n5340 VDD.n5338 1.49065
R4357 VDD.n5336 VDD.n5334 1.49065
R4358 VDD.n5332 VDD.n5330 1.49065
R4359 VDD.n5328 VDD.n5326 1.49065
R4360 VDD.n5324 VDD.n5322 1.49065
R4361 VDD.n5320 VDD.n5318 1.49065
R4362 VDD.n5316 VDD.n5314 1.49065
R4363 VDD.n5312 VDD.n5310 1.49065
R4364 VDD.n5308 VDD.n5306 1.49065
R4365 VDD.n5304 VDD.n5302 1.49065
R4366 VDD.n5300 VDD.n5298 1.49065
R4367 VDD.n5296 VDD.n5294 1.49065
R4368 VDD.n5292 VDD.n5290 1.49065
R4369 VDD.n5288 VDD.n5286 1.49065
R4370 VDD.n5284 VDD.n5282 1.49065
R4371 VDD.n13 VDD.n11 1.49065
R4372 VDD.n17 VDD.n15 1.49065
R4373 VDD.n21 VDD.n19 1.49065
R4374 VDD.n25 VDD.n23 1.49065
R4375 VDD.n29 VDD.n27 1.49065
R4376 VDD.n33 VDD.n31 1.49065
R4377 VDD.n37 VDD.n35 1.49065
R4378 VDD.n41 VDD.n39 1.49065
R4379 VDD.n45 VDD.n43 1.49065
R4380 VDD.n49 VDD.n47 1.49065
R4381 VDD.n53 VDD.n51 1.49065
R4382 VDD.n57 VDD.n55 1.49065
R4383 VDD.n61 VDD.n59 1.49065
R4384 VDD.n65 VDD.n63 1.49065
R4385 VDD.n69 VDD.n67 1.49065
R4386 VDD.n3416 VDD.n3415 1.4691
R4387 VDD.n3439 VDD.n3437 1.4691
R4388 VDD.n3611 VDD.n3609 1.4691
R4389 VDD.n3778 VDD.n3777 1.4691
R4390 VDD.n3800 VDD.n3798 1.4691
R4391 VDD.n3968 VDD.n3966 1.4691
R4392 VDD.n4129 VDD.n4128 1.4691
R4393 VDD.n4149 VDD.n4148 1.4691
R4394 VDD.n4299 VDD.n4298 1.4691
R4395 VDD.n4397 VDD.t27 1.4691
R4396 VDD.n4450 VDD.n4449 1.4691
R4397 VDD.n4473 VDD.n4471 1.4691
R4398 VDD.n4542 VDD.t50 1.4691
R4399 VDD.n4643 VDD.n4641 1.4691
R4400 VDD.n4803 VDD.n4802 1.4691
R4401 VDD.n4829 VDD.n4827 1.4691
R4402 VDD.n5001 VDD.n4999 1.4691
R4403 VDD.n5157 VDD.n5156 1.4691
R4404 VDD.n6783 VDD.n6782 1.43601
R4405 VDD.n941 VDD.n940 1.43109
R4406 VDD.n1519 VDD.n1518 1.4204
R4407 VDD.n3 VDD.n1 1.4204
R4408 VDD.n5 VDD.n3 1.4204
R4409 VDD.n7 VDD.n5 1.4204
R4410 VDD.n9 VDD.n7 1.4204
R4411 VDD.n89 VDD.n87 1.4204
R4412 VDD.n85 VDD.n84 1.41423
R4413 VDD.n1796 VDD.n1795 1.40363
R4414 VDD.n1521 VDD.n1519 1.39758
R4415 VDD.n180 VDD.n179 1.39686
R4416 VDD.n223 VDD.n222 1.39686
R4417 VDD.n261 VDD.n169 1.39686
R4418 VDD.n1193 VDD.n1191 1.39537
R4419 VDD.n1205 VDD.n1203 1.39537
R4420 VDD.n1203 VDD.n1201 1.39537
R4421 VDD.n1201 VDD.n1199 1.39537
R4422 VDD.n1199 VDD.n1197 1.39537
R4423 VDD.n1197 VDD.n1195 1.39537
R4424 VDD.n1213 VDD.n1211 1.39537
R4425 VDD.n1215 VDD.n1213 1.39537
R4426 VDD.n1217 VDD.n1215 1.39537
R4427 VDD.n1219 VDD.n1217 1.39537
R4428 VDD.n1221 VDD.n1219 1.39537
R4429 VDD.n1319 VDD.n1317 1.39537
R4430 VDD.n1294 VDD.n1292 1.39537
R4431 VDD.n1289 VDD.n1287 1.39537
R4432 VDD.n1746 VDD.n1744 1.39537
R4433 VDD.n1751 VDD.n1749 1.39537
R4434 VDD.n1789 VDD.n1787 1.39537
R4435 VDD.n1625 VDD.n1623 1.39537
R4436 VDD.n1620 VDD.n1618 1.39537
R4437 VDD.n1583 VDD.n1581 1.39537
R4438 VDD.n1578 VDD.n1576 1.39537
R4439 VDD.n1477 VDD.n1475 1.39537
R4440 VDD.n1509 VDD.n1507 1.39537
R4441 VDD.n1514 VDD.n1512 1.39537
R4442 VDD.n1523 VDD.n1521 1.39537
R4443 VDD.n1257 VDD.n1255 1.35435
R4444 VDD.n815 VDD.n814 1.35205
R4445 VDD.n727 VDD.n726 1.35205
R4446 VDD.n639 VDD.n638 1.35205
R4447 VDD.n551 VDD.n550 1.35205
R4448 VDD.n463 VDD.n462 1.35205
R4449 VDD.n6364 VDD.n6359 1.33781
R4450 VDD.n6259 VDD.n6254 1.33781
R4451 VDD.n321 VDD.n320 1.31929
R4452 VDD.n366 VDD.n365 1.31929
R4453 VDD.n1655 VDD.n1653 1.31332
R4454 VDD.n1649 VDD.n1647 1.31332
R4455 VDD.n1643 VDD.n1641 1.31332
R4456 VDD.n1637 VDD.n1635 1.31332
R4457 VDD.n1631 VDD.n1629 1.31332
R4458 VDD.n6378 VDD.n6377 1.2996
R4459 VDD.n6272 VDD.n6271 1.2996
R4460 VDD.n3591 VDD.n3587 1.28552
R4461 VDD.n3630 VDD.n3629 1.28552
R4462 VDD.n3650 VDD.t17 1.28552
R4463 VDD.n3781 VDD.n3780 1.28552
R4464 VDD.n3951 VDD.n3947 1.28552
R4465 VDD.t11 VDD.n3968 1.28552
R4466 VDD.n3994 VDD.n3993 1.28552
R4467 VDD.n4131 VDD.n4130 1.28552
R4468 VDD.t105 VDD.n4242 1.28552
R4469 VDD.n4261 VDD.t13 1.28552
R4470 VDD.n4279 VDD.n4276 1.28552
R4471 VDD.n4322 VDD.n4321 1.28552
R4472 VDD.n4453 VDD.n4452 1.28552
R4473 VDD.t50 VDD.n4537 1.28552
R4474 VDD.n4667 VDD.n4666 1.28552
R4475 VDD.n4978 VDD.n4974 1.28552
R4476 VDD.n5023 VDD.n5022 1.28552
R4477 VDD.n5263 VDD.n5158 1.28552
R4478 VDD.n6698 VDD.n6697 1.28539
R4479 VDD.n3473 VDD.n3472 1.2805
R4480 VDD.n3511 VDD.n3510 1.2805
R4481 VDD.n3574 VDD.n3561 1.2805
R4482 VDD.n3563 VDD.n3562 1.2805
R4483 VDD.n3657 VDD.n3656 1.2805
R4484 VDD.n3825 VDD.n3824 1.2805
R4485 VDD.n3837 VDD.n3836 1.2805
R4486 VDD.n3893 VDD.n3890 1.2805
R4487 VDD.n3933 VDD.n3920 1.2805
R4488 VDD.n3922 VDD.n3921 1.2805
R4489 VDD.n3977 VDD.n3976 1.2805
R4490 VDD.n4020 VDD.n4010 1.2805
R4491 VDD.n4135 VDD.n4133 1.2805
R4492 VDD.n4184 VDD.n4183 1.2805
R4493 VDD.n4200 VDD.n4199 1.2805
R4494 VDD.n4266 VDD.n4255 1.2805
R4495 VDD.n4257 VDD.n4256 1.2805
R4496 VDD.n4484 VDD.n4483 1.2805
R4497 VDD.n4501 VDD.n4500 1.2805
R4498 VDD.n4500 VDD.n4490 1.2805
R4499 VDD.n4512 VDD.n4511 1.2805
R4500 VDD.n4602 VDD.n4601 1.2805
R4501 VDD.n4793 VDD.n4792 1.2805
R4502 VDD.n4809 VDD.n4808 1.2805
R4503 VDD.n4864 VDD.n4863 1.2805
R4504 VDD.n4876 VDD.n4875 1.2805
R4505 VDD.n4957 VDD.n4947 1.2805
R4506 VDD.n4959 VDD.n4958 1.2805
R4507 VDD.n6786 VDD.n6783 1.27651
R4508 VDD.n1473 VDD.n1472 1.27229
R4509 VDD.n6498 VDD.n6485 1.26018
R4510 VDD.n1320 VDD.n1319 1.25178
R4511 VDD.n1452 VDD.n1450 1.23127
R4512 VDD.n1457 VDD.n1455 1.23127
R4513 VDD.n1462 VDD.n1460 1.23127
R4514 VDD.n1467 VDD.n1465 1.23127
R4515 VDD.n1472 VDD.n1470 1.23127
R4516 VDD.n2830 VDD.n2828 1.22558
R4517 VDD.n2826 VDD.n2824 1.22558
R4518 VDD.n2823 VDD.n2821 1.22558
R4519 VDD.n2820 VDD.n2818 1.22558
R4520 VDD.n2817 VDD.n2815 1.22558
R4521 VDD.n2814 VDD.n2812 1.22558
R4522 VDD.n2811 VDD.n2809 1.22558
R4523 VDD.n2808 VDD.n2806 1.22558
R4524 VDD.n2805 VDD.n2803 1.22558
R4525 VDD.n2802 VDD.n2800 1.22558
R4526 VDD.n2799 VDD.n2797 1.22558
R4527 VDD.n2796 VDD.n2794 1.22558
R4528 VDD.n2793 VDD.n2791 1.22558
R4529 VDD.n2790 VDD.n2788 1.22558
R4530 VDD.n1021 VDD.n1020 1.22558
R4531 VDD.n1024 VDD.n1023 1.22558
R4532 VDD.n1027 VDD.n1026 1.22558
R4533 VDD.n1030 VDD.n1029 1.22558
R4534 VDD.n1033 VDD.n1032 1.22558
R4535 VDD.n1036 VDD.n1035 1.22558
R4536 VDD.n1039 VDD.n1038 1.22558
R4537 VDD.n1042 VDD.n1041 1.22558
R4538 VDD.n1045 VDD.n1044 1.22558
R4539 VDD.n1048 VDD.n1047 1.22558
R4540 VDD.n1051 VDD.n1050 1.22558
R4541 VDD.n1054 VDD.n1053 1.22558
R4542 VDD.n1058 VDD.n1056 1.22558
R4543 VDD.n1062 VDD.n1060 1.22558
R4544 VDD.n1066 VDD.n1064 1.22558
R4545 VDD.n1070 VDD.n1068 1.22558
R4546 VDD.n1074 VDD.n1072 1.22558
R4547 VDD.n1078 VDD.n1076 1.22558
R4548 VDD.n863 VDD.n862 1.19305
R4549 VDD.n775 VDD.n774 1.19305
R4550 VDD.n687 VDD.n686 1.19305
R4551 VDD.n599 VDD.n598 1.19305
R4552 VDD.n511 VDD.n510 1.19305
R4553 VDD.n423 VDD.n422 1.19305
R4554 VDD.n1792 VDD.n1790 1.19024
R4555 VDD.n6370 VDD.n6367 1.18498
R4556 VDD.n6264 VDD.n6261 1.18498
R4557 VDD.n85 VDD.n81 1.18498
R4558 VDD.n1285 VDD.n1282 1.14922
R4559 VDD.n1280 VDD.n1277 1.14922
R4560 VDD.n1275 VDD.n1272 1.14922
R4561 VDD.n1270 VDD.n1267 1.14922
R4562 VDD.n1265 VDD.n1262 1.14922
R4563 VDD.n1260 VDD.n1257 1.14922
R4564 VDD.n6370 VDD.n6369 1.14677
R4565 VDD.n6264 VDD.n6263 1.14677
R4566 VDD.n6252 VDD.n6080 1.14433
R4567 VDD.n6250 VDD.n6087 1.14433
R4568 VDD.n6248 VDD.n6094 1.14433
R4569 VDD.n6246 VDD.n6101 1.14433
R4570 VDD.n6244 VDD.n6108 1.14433
R4571 VDD.n6242 VDD.n6115 1.14433
R4572 VDD.n6240 VDD.n6122 1.14433
R4573 VDD.n6238 VDD.n6129 1.14433
R4574 VDD.n6236 VDD.n6136 1.14433
R4575 VDD.n6234 VDD.n6143 1.14433
R4576 VDD.n6232 VDD.n6150 1.14433
R4577 VDD.n6230 VDD.n6157 1.14433
R4578 VDD.n6228 VDD.n6164 1.14433
R4579 VDD.n6226 VDD.n6171 1.14433
R4580 VDD.n6224 VDD.n6178 1.14433
R4581 VDD.n6222 VDD.n6185 1.14433
R4582 VDD.n6220 VDD.n6192 1.14433
R4583 VDD.n6218 VDD.n6199 1.14433
R4584 VDD.n6216 VDD.n6206 1.14433
R4585 VDD.n6214 VDD.n6213 1.14433
R4586 VDD.n6073 VDD.n5901 1.14433
R4587 VDD.n6071 VDD.n5908 1.14433
R4588 VDD.n6069 VDD.n5915 1.14433
R4589 VDD.n6067 VDD.n5922 1.14433
R4590 VDD.n6065 VDD.n5929 1.14433
R4591 VDD.n6063 VDD.n5936 1.14433
R4592 VDD.n6061 VDD.n5943 1.14433
R4593 VDD.n6059 VDD.n5950 1.14433
R4594 VDD.n6057 VDD.n5957 1.14433
R4595 VDD.n6055 VDD.n5964 1.14433
R4596 VDD.n6053 VDD.n5971 1.14433
R4597 VDD.n6051 VDD.n5978 1.14433
R4598 VDD.n6049 VDD.n5985 1.14433
R4599 VDD.n6047 VDD.n5992 1.14433
R4600 VDD.n6045 VDD.n5999 1.14433
R4601 VDD.n6043 VDD.n6006 1.14433
R4602 VDD.n6041 VDD.n6013 1.14433
R4603 VDD.n6039 VDD.n6020 1.14433
R4604 VDD.n6037 VDD.n6027 1.14433
R4605 VDD.n6035 VDD.n6034 1.14433
R4606 VDD.n5894 VDD.n5722 1.14433
R4607 VDD.n5892 VDD.n5729 1.14433
R4608 VDD.n5890 VDD.n5736 1.14433
R4609 VDD.n5888 VDD.n5743 1.14433
R4610 VDD.n5886 VDD.n5750 1.14433
R4611 VDD.n5884 VDD.n5757 1.14433
R4612 VDD.n5882 VDD.n5764 1.14433
R4613 VDD.n5880 VDD.n5771 1.14433
R4614 VDD.n5878 VDD.n5778 1.14433
R4615 VDD.n5876 VDD.n5785 1.14433
R4616 VDD.n5874 VDD.n5792 1.14433
R4617 VDD.n5872 VDD.n5799 1.14433
R4618 VDD.n5870 VDD.n5806 1.14433
R4619 VDD.n5868 VDD.n5813 1.14433
R4620 VDD.n5866 VDD.n5820 1.14433
R4621 VDD.n5864 VDD.n5827 1.14433
R4622 VDD.n5862 VDD.n5834 1.14433
R4623 VDD.n5860 VDD.n5841 1.14433
R4624 VDD.n5858 VDD.n5848 1.14433
R4625 VDD.n5856 VDD.n5855 1.14433
R4626 VDD.n5715 VDD.n5543 1.14433
R4627 VDD.n5713 VDD.n5550 1.14433
R4628 VDD.n5711 VDD.n5557 1.14433
R4629 VDD.n5709 VDD.n5564 1.14433
R4630 VDD.n5707 VDD.n5571 1.14433
R4631 VDD.n5705 VDD.n5578 1.14433
R4632 VDD.n5703 VDD.n5585 1.14433
R4633 VDD.n5701 VDD.n5592 1.14433
R4634 VDD.n5699 VDD.n5599 1.14433
R4635 VDD.n5697 VDD.n5606 1.14433
R4636 VDD.n5695 VDD.n5613 1.14433
R4637 VDD.n5693 VDD.n5620 1.14433
R4638 VDD.n5691 VDD.n5627 1.14433
R4639 VDD.n5689 VDD.n5634 1.14433
R4640 VDD.n5687 VDD.n5641 1.14433
R4641 VDD.n5685 VDD.n5648 1.14433
R4642 VDD.n5683 VDD.n5655 1.14433
R4643 VDD.n5681 VDD.n5662 1.14433
R4644 VDD.n5679 VDD.n5669 1.14433
R4645 VDD.n5677 VDD.n5676 1.14433
R4646 VDD.n5536 VDD.n5364 1.14433
R4647 VDD.n5534 VDD.n5371 1.14433
R4648 VDD.n5532 VDD.n5378 1.14433
R4649 VDD.n5530 VDD.n5385 1.14433
R4650 VDD.n5528 VDD.n5392 1.14433
R4651 VDD.n5526 VDD.n5399 1.14433
R4652 VDD.n5524 VDD.n5406 1.14433
R4653 VDD.n5522 VDD.n5413 1.14433
R4654 VDD.n5520 VDD.n5420 1.14433
R4655 VDD.n5518 VDD.n5427 1.14433
R4656 VDD.n5516 VDD.n5434 1.14433
R4657 VDD.n5514 VDD.n5441 1.14433
R4658 VDD.n5512 VDD.n5448 1.14433
R4659 VDD.n5510 VDD.n5455 1.14433
R4660 VDD.n5508 VDD.n5462 1.14433
R4661 VDD.n5506 VDD.n5469 1.14433
R4662 VDD.n5504 VDD.n5476 1.14433
R4663 VDD.n5502 VDD.n5483 1.14433
R4664 VDD.n5500 VDD.n5490 1.14433
R4665 VDD.n5498 VDD.n5497 1.14433
R4666 VDD.n2691 VDD.n2519 1.14433
R4667 VDD.n2689 VDD.n2526 1.14433
R4668 VDD.n2687 VDD.n2533 1.14433
R4669 VDD.n2685 VDD.n2540 1.14433
R4670 VDD.n2683 VDD.n2547 1.14433
R4671 VDD.n2681 VDD.n2554 1.14433
R4672 VDD.n2679 VDD.n2561 1.14433
R4673 VDD.n2677 VDD.n2568 1.14433
R4674 VDD.n2675 VDD.n2575 1.14433
R4675 VDD.n2673 VDD.n2582 1.14433
R4676 VDD.n2671 VDD.n2589 1.14433
R4677 VDD.n2669 VDD.n2596 1.14433
R4678 VDD.n2667 VDD.n2603 1.14433
R4679 VDD.n2665 VDD.n2610 1.14433
R4680 VDD.n2663 VDD.n2617 1.14433
R4681 VDD.n2661 VDD.n2624 1.14433
R4682 VDD.n2659 VDD.n2631 1.14433
R4683 VDD.n2657 VDD.n2638 1.14433
R4684 VDD.n2655 VDD.n2645 1.14433
R4685 VDD.n2653 VDD.n2652 1.14433
R4686 VDD.n2512 VDD.n2340 1.14433
R4687 VDD.n2510 VDD.n2347 1.14433
R4688 VDD.n2508 VDD.n2354 1.14433
R4689 VDD.n2506 VDD.n2361 1.14433
R4690 VDD.n2504 VDD.n2368 1.14433
R4691 VDD.n2502 VDD.n2375 1.14433
R4692 VDD.n2500 VDD.n2382 1.14433
R4693 VDD.n2498 VDD.n2389 1.14433
R4694 VDD.n2496 VDD.n2396 1.14433
R4695 VDD.n2494 VDD.n2403 1.14433
R4696 VDD.n2492 VDD.n2410 1.14433
R4697 VDD.n2490 VDD.n2417 1.14433
R4698 VDD.n2488 VDD.n2424 1.14433
R4699 VDD.n2486 VDD.n2431 1.14433
R4700 VDD.n2484 VDD.n2438 1.14433
R4701 VDD.n2482 VDD.n2445 1.14433
R4702 VDD.n2480 VDD.n2452 1.14433
R4703 VDD.n2478 VDD.n2459 1.14433
R4704 VDD.n2476 VDD.n2466 1.14433
R4705 VDD.n2474 VDD.n2473 1.14433
R4706 VDD.n2333 VDD.n2161 1.14433
R4707 VDD.n2331 VDD.n2168 1.14433
R4708 VDD.n2329 VDD.n2175 1.14433
R4709 VDD.n2327 VDD.n2182 1.14433
R4710 VDD.n2325 VDD.n2189 1.14433
R4711 VDD.n2323 VDD.n2196 1.14433
R4712 VDD.n2321 VDD.n2203 1.14433
R4713 VDD.n2319 VDD.n2210 1.14433
R4714 VDD.n2317 VDD.n2217 1.14433
R4715 VDD.n2315 VDD.n2224 1.14433
R4716 VDD.n2313 VDD.n2231 1.14433
R4717 VDD.n2311 VDD.n2238 1.14433
R4718 VDD.n2309 VDD.n2245 1.14433
R4719 VDD.n2307 VDD.n2252 1.14433
R4720 VDD.n2305 VDD.n2259 1.14433
R4721 VDD.n2303 VDD.n2266 1.14433
R4722 VDD.n2301 VDD.n2273 1.14433
R4723 VDD.n2299 VDD.n2280 1.14433
R4724 VDD.n2297 VDD.n2287 1.14433
R4725 VDD.n2295 VDD.n2294 1.14433
R4726 VDD.n2154 VDD.n1982 1.14433
R4727 VDD.n2152 VDD.n1989 1.14433
R4728 VDD.n2150 VDD.n1996 1.14433
R4729 VDD.n2148 VDD.n2003 1.14433
R4730 VDD.n2146 VDD.n2010 1.14433
R4731 VDD.n2144 VDD.n2017 1.14433
R4732 VDD.n2142 VDD.n2024 1.14433
R4733 VDD.n2140 VDD.n2031 1.14433
R4734 VDD.n2138 VDD.n2038 1.14433
R4735 VDD.n2136 VDD.n2045 1.14433
R4736 VDD.n2134 VDD.n2052 1.14433
R4737 VDD.n2132 VDD.n2059 1.14433
R4738 VDD.n2130 VDD.n2066 1.14433
R4739 VDD.n2128 VDD.n2073 1.14433
R4740 VDD.n2126 VDD.n2080 1.14433
R4741 VDD.n2124 VDD.n2087 1.14433
R4742 VDD.n2122 VDD.n2094 1.14433
R4743 VDD.n2120 VDD.n2101 1.14433
R4744 VDD.n2118 VDD.n2108 1.14433
R4745 VDD.n2116 VDD.n2115 1.14433
R4746 VDD.n1975 VDD.n1803 1.14433
R4747 VDD.n1973 VDD.n1810 1.14433
R4748 VDD.n1971 VDD.n1817 1.14433
R4749 VDD.n1969 VDD.n1824 1.14433
R4750 VDD.n1967 VDD.n1831 1.14433
R4751 VDD.n1965 VDD.n1838 1.14433
R4752 VDD.n1963 VDD.n1845 1.14433
R4753 VDD.n1961 VDD.n1852 1.14433
R4754 VDD.n1959 VDD.n1859 1.14433
R4755 VDD.n1957 VDD.n1866 1.14433
R4756 VDD.n1955 VDD.n1873 1.14433
R4757 VDD.n1953 VDD.n1880 1.14433
R4758 VDD.n1951 VDD.n1887 1.14433
R4759 VDD.n1949 VDD.n1894 1.14433
R4760 VDD.n1947 VDD.n1901 1.14433
R4761 VDD.n1945 VDD.n1908 1.14433
R4762 VDD.n1943 VDD.n1915 1.14433
R4763 VDD.n1941 VDD.n1922 1.14433
R4764 VDD.n1939 VDD.n1929 1.14433
R4765 VDD.n1937 VDD.n1936 1.14433
R4766 VDD.n946 VDD.n945 1.12991
R4767 VDD.n109 VDD.n108 1.12832
R4768 VDD.n6697 VDD.n6505 1.11501
R4769 VDD.n375 VDD.n374 1.11354
R4770 VDD.n5350 VDD.n5348 1.10856
R4771 VDD.n5346 VDD.n5344 1.10856
R4772 VDD.n5342 VDD.n5340 1.10856
R4773 VDD.n5338 VDD.n5336 1.10856
R4774 VDD.n5334 VDD.n5332 1.10856
R4775 VDD.n5330 VDD.n5328 1.10856
R4776 VDD.n5326 VDD.n5324 1.10856
R4777 VDD.n5322 VDD.n5320 1.10856
R4778 VDD.n5318 VDD.n5316 1.10856
R4779 VDD.n5314 VDD.n5312 1.10856
R4780 VDD.n5310 VDD.n5308 1.10856
R4781 VDD.n5306 VDD.n5304 1.10856
R4782 VDD.n5302 VDD.n5300 1.10856
R4783 VDD.n5298 VDD.n5296 1.10856
R4784 VDD.n5294 VDD.n5292 1.10856
R4785 VDD.n5290 VDD.n5288 1.10856
R4786 VDD.n5286 VDD.n5284 1.10856
R4787 VDD.n15 VDD.n13 1.10856
R4788 VDD.n19 VDD.n17 1.10856
R4789 VDD.n23 VDD.n21 1.10856
R4790 VDD.n27 VDD.n25 1.10856
R4791 VDD.n31 VDD.n29 1.10856
R4792 VDD.n35 VDD.n33 1.10856
R4793 VDD.n39 VDD.n37 1.10856
R4794 VDD.n43 VDD.n41 1.10856
R4795 VDD.n47 VDD.n45 1.10856
R4796 VDD.n51 VDD.n49 1.10856
R4797 VDD.n55 VDD.n53 1.10856
R4798 VDD.n59 VDD.n57 1.10856
R4799 VDD.n63 VDD.n61 1.10856
R4800 VDD.n67 VDD.n65 1.10856
R4801 VDD.n3396 VDD.n3395 1.10195
R4802 VDD.n3419 VDD.t61 1.10195
R4803 VDD.n3459 VDD.n3457 1.10195
R4804 VDD.n3590 VDD.n3588 1.10195
R4805 VDD.n3758 VDD.n3757 1.10195
R4806 VDD.n3821 VDD.n3819 1.10195
R4807 VDD.n3950 VDD.n3948 1.10195
R4808 VDD.n4111 VDD.n4110 1.10195
R4809 VDD.n4170 VDD.n4169 1.10195
R4810 VDD.n4278 VDD.n4277 1.10195
R4811 VDD.n4432 VDD.n4431 1.10195
R4812 VDD.n4497 VDD.n4495 1.10195
R4813 VDD.n4621 VDD.t115 1.10195
R4814 VDD.n4620 VDD.n4618 1.10195
R4815 VDD.n4780 VDD.n4779 1.10195
R4816 VDD.n4852 VDD.n4850 1.10195
R4817 VDD.n4977 VDD.n4975 1.10195
R4818 VDD.n5134 VDD.n5133 1.10195
R4819 VDD.n176 VDD.n175 1.08656
R4820 VDD.n228 VDD.n227 1.08656
R4821 VDD.n166 VDD.n165 1.08656
R4822 VDD.n1714 VDD.n1711 1.06717
R4823 VDD.n1719 VDD.n1716 1.06717
R4824 VDD.n1724 VDD.n1721 1.06717
R4825 VDD.n1730 VDD.n1726 1.06717
R4826 VDD.n1736 VDD.n1732 1.06717
R4827 VDD.n1742 VDD.n1738 1.06717
R4828 VDD.n1314 VDD.n1312 1.04665
R4829 VDD.n1309 VDD.n1307 1.04665
R4830 VDD.n1304 VDD.n1302 1.04665
R4831 VDD.n1299 VDD.n1297 1.04665
R4832 VDD.n810 VDD.n809 1.03404
R4833 VDD.n722 VDD.n721 1.03404
R4834 VDD.n634 VDD.n633 1.03404
R4835 VDD.n546 VDD.n545 1.03404
R4836 VDD.n458 VDD.n457 1.03404
R4837 VDD.n6378 VDD.n6375 1.03214
R4838 VDD.n6272 VDD.n6269 1.03214
R4839 VDD.n1623 VDD.n1621 1.02614
R4840 VDD.n316 VDD.n315 1.00898
R4841 VDD.n6364 VDD.n6363 0.993933
R4842 VDD.n6259 VDD.n6258 0.993933
R4843 VDD.n1480 VDD.n1477 0.985115
R4844 VDD.n1485 VDD.n1482 0.985115
R4845 VDD.n1490 VDD.n1487 0.985115
R4846 VDD.n1495 VDD.n1492 0.985115
R4847 VDD.n1500 VDD.n1497 0.985115
R4848 VDD.n1505 VDD.n1502 0.985115
R4849 VDD.n2833 VDD.n2832 0.972117
R4850 VDD.n3045 VDD.n3043 0.9605
R4851 VDD.n3016 VDD.n3006 0.9605
R4852 VDD.n3666 VDD.n3665 0.9605
R4853 VDD.n3681 VDD.n3680 0.9605
R4854 VDD.n3743 VDD.n3733 0.9605
R4855 VDD.n3745 VDD.n3743 0.9605
R4856 VDD.n3830 VDD.n3829 0.9605
R4857 VDD.n3853 VDD.n3852 0.9605
R4858 VDD.n3983 VDD.n3982 0.9605
R4859 VDD.n4043 VDD.n4042 0.9605
R4860 VDD.n4096 VDD.n4088 0.9605
R4861 VDD.n4098 VDD.n4096 0.9605
R4862 VDD.n4282 VDD.n4273 0.9605
R4863 VDD.n4333 VDD.n4332 0.9605
R4864 VDD.n4348 VDD.n4345 0.9605
R4865 VDD.n4418 VDD.n4410 0.9605
R4866 VDD.n4420 VDD.n4418 0.9605
R4867 VDD.n4631 VDD.n4630 0.9605
R4868 VDD.n4649 VDD.n4646 0.9605
R4869 VDD.n4654 VDD.n4653 0.9605
R4870 VDD.n4711 VDD.n4710 0.9605
R4871 VDD.n4710 VDD.n4700 0.9605
R4872 VDD.n4768 VDD.n4758 0.9605
R4873 VDD.n4786 VDD.n4775 0.9605
R4874 VDD.n4792 VDD.n4791 0.9605
R4875 VDD.n4809 VDD.n4798 0.9605
R4876 VDD.n4835 VDD.n4821 0.9605
R4877 VDD.n4942 VDD.n4941 0.9605
R4878 VDD.n4960 VDD.n4957 0.9605
R4879 VDD.n5026 VDD.n5025 0.9605
R4880 VDD.n5065 VDD.n5064 0.9605
R4881 VDD.n5064 VDD.n5054 0.9605
R4882 VDD.n5118 VDD.n5117 0.9605
R4883 VDD.n1579 VDD.n1578 0.94409
R4884 VDD.n1512 VDD.n1510 0.94409
R4885 VDD.n1795 VDD.n1208 0.91841
R4886 VDD.n3399 VDD.n3398 0.918374
R4887 VDD.t45 VDD.n3507 0.918374
R4888 VDD.n3571 VDD.n3567 0.918374
R4889 VDD.n3654 VDD.n3653 0.918374
R4890 VDD.n3761 VDD.n3760 0.918374
R4891 VDD.n3930 VDD.n3926 0.918374
R4892 VDD.n4018 VDD.n4017 0.918374
R4893 VDD.n4113 VDD.n4112 0.918374
R4894 VDD.n4263 VDD.n4260 0.918374
R4895 VDD.n4343 VDD.n4342 0.918374
R4896 VDD.t78 VDD.n4359 0.918374
R4897 VDD.n4434 VDD.n4433 0.918374
R4898 VDD.n4597 VDD.n4593 0.918374
R4899 VDD.n4666 VDD.t93 0.918374
R4900 VDD.t93 VDD.n4664 0.918374
R4901 VDD.n4689 VDD.n4688 0.918374
R4902 VDD.n4783 VDD.n4782 0.918374
R4903 VDD.n4955 VDD.n4951 0.918374
R4904 VDD.n5038 VDD.t117 0.918374
R4905 VDD.n5042 VDD.n5041 0.918374
R4906 VDD.n5136 VDD.n5135 0.918374
R4907 VDD.n6790 VDD.n6789 0.917515
R4908 VDD.n1757 VDD.n1755 0.903064
R4909 VDD.n1763 VDD.n1761 0.903064
R4910 VDD.n1769 VDD.n1767 0.903064
R4911 VDD.n1775 VDD.n1773 0.903064
R4912 VDD.n1781 VDD.n1779 0.903064
R4913 VDD.n1787 VDD.n1785 0.903064
R4914 VDD.n6384 VDD.n6383 0.879306
R4915 VDD.n6278 VDD.n6277 0.879306
R4916 VDD.n5353 VDD.n5352 0.879306
R4917 VDD.n780 VDD.n779 0.875034
R4918 VDD.n692 VDD.n691 0.875034
R4919 VDD.n604 VDD.n603 0.875034
R4920 VDD.n516 VDD.n515 0.875034
R4921 VDD.n428 VDD.n427 0.875034
R4922 VDD.n1206 VDD.n1193 0.862038
R4923 VDD.n1290 VDD.n1289 0.862038
R4924 VDD.n1315 VDD.n1314 0.841526
R4925 VDD.n6356 VDD.n6355 0.841097
R4926 VDD.n1017 VDD.n1016 0.828735
R4927 VDD.n1515 VDD.n1514 0.821013
R4928 VDD.n3048 VDD.n3047 0.819831
R4929 VDD.n1747 VDD.n1746 0.779987
R4930 VDD.n233 VDD.n232 0.776258
R4931 VDD.n258 VDD.n257 0.776258
R4932 VDD.n90 VDD.n9 0.773094
R4933 VDD.n1660 VDD.n1659 0.759474
R4934 VDD.n1618 VDD.n1616 0.738962
R4935 VDD.n1612 VDD.n1610 0.738962
R4936 VDD.n1606 VDD.n1604 0.738962
R4937 VDD.n1600 VDD.n1598 0.738962
R4938 VDD.n1594 VDD.n1592 0.738962
R4939 VDD.n1588 VDD.n1586 0.738962
R4940 VDD.n3011 VDD.n3010 0.734799
R4941 VDD.n3480 VDD.n3478 0.734799
R4942 VDD.n3570 VDD.n3568 0.734799
R4943 VDD.n3738 VDD.n3737 0.734799
R4944 VDD.n3844 VDD.n3842 0.734799
R4945 VDD.n3929 VDD.n3927 0.734799
R4946 VDD.n4092 VDD.n4091 0.734799
R4947 VDD.n4150 VDD.t133 0.734799
R4948 VDD.n4189 VDD.n4188 0.734799
R4949 VDD.n4262 VDD.n4261 0.734799
R4950 VDD.n4414 VDD.n4413 0.734799
R4951 VDD.n4519 VDD.n4517 0.734799
R4952 VDD.n4596 VDD.n4594 0.734799
R4953 VDD.n4763 VDD.n4762 0.734799
R4954 VDD.n4806 VDD.t2 0.734799
R4955 VDD.n4871 VDD.n4869 0.734799
R4956 VDD.n4954 VDD.n4952 0.734799
R4957 VDD.n5113 VDD.n5112 0.734799
R4958 VDD.n2697 VDD.n2696 0.731929
R4959 VDD.n6508 VDD.n6507 0.731929
R4960 VDD.n6510 VDD.n6509 0.731929
R4961 VDD.n6512 VDD.n6511 0.731929
R4962 VDD.n6514 VDD.n6513 0.731929
R4963 VDD.n6516 VDD.n6515 0.731929
R4964 VDD.n6518 VDD.n6517 0.731929
R4965 VDD.n6520 VDD.n6519 0.731929
R4966 VDD.n6522 VDD.n6521 0.731929
R4967 VDD.n6524 VDD.n6523 0.731929
R4968 VDD.n6526 VDD.n6525 0.731929
R4969 VDD.n6528 VDD.n6527 0.731929
R4970 VDD.n6530 VDD.n6529 0.731929
R4971 VDD.n6532 VDD.n6531 0.731929
R4972 VDD.n6534 VDD.n6533 0.731929
R4973 VDD.n6536 VDD.n6535 0.731929
R4974 VDD.n6538 VDD.n6537 0.731929
R4975 VDD.n6540 VDD.n6539 0.731929
R4976 VDD.n6542 VDD.n6541 0.731929
R4977 VDD.n6544 VDD.n6543 0.731929
R4978 VDD.n6546 VDD.n6545 0.731929
R4979 VDD.n6548 VDD.n6547 0.731929
R4980 VDD.n6550 VDD.n6549 0.731929
R4981 VDD.n6552 VDD.n6551 0.731929
R4982 VDD.n6554 VDD.n6553 0.731929
R4983 VDD.n6556 VDD.n6555 0.731929
R4984 VDD.n6558 VDD.n6557 0.731929
R4985 VDD.n6560 VDD.n6559 0.731929
R4986 VDD.n6562 VDD.n6561 0.731929
R4987 VDD.n6564 VDD.n6563 0.731929
R4988 VDD.n6566 VDD.n6565 0.731929
R4989 VDD.n6568 VDD.n6567 0.731929
R4990 VDD.n6570 VDD.n6569 0.731929
R4991 VDD.n6572 VDD.n6571 0.731929
R4992 VDD.n6575 VDD.n6574 0.731929
R4993 VDD.n6579 VDD.n6577 0.731929
R4994 VDD.n6583 VDD.n6581 0.731929
R4995 VDD.n6587 VDD.n6585 0.731929
R4996 VDD.n6591 VDD.n6589 0.731929
R4997 VDD.n6595 VDD.n6593 0.731929
R4998 VDD.n6599 VDD.n6597 0.731929
R4999 VDD.n6603 VDD.n6601 0.731929
R5000 VDD.n6607 VDD.n6605 0.731929
R5001 VDD.n6611 VDD.n6609 0.731929
R5002 VDD.n6615 VDD.n6613 0.731929
R5003 VDD.n6619 VDD.n6617 0.731929
R5004 VDD.n6693 VDD.n6691 0.731929
R5005 VDD.n6689 VDD.n6687 0.731929
R5006 VDD.n6685 VDD.n6683 0.731929
R5007 VDD.n6681 VDD.n6679 0.731929
R5008 VDD.n6677 VDD.n6675 0.731929
R5009 VDD.n6673 VDD.n6671 0.731929
R5010 VDD.n6669 VDD.n6667 0.731929
R5011 VDD.n6665 VDD.n6663 0.731929
R5012 VDD.n6661 VDD.n6659 0.731929
R5013 VDD.n6657 VDD.n6655 0.731929
R5014 VDD.n6653 VDD.n6651 0.731929
R5015 VDD.n6650 VDD.n6649 0.731929
R5016 VDD.n6648 VDD.n6647 0.731929
R5017 VDD.n6646 VDD.n6645 0.731929
R5018 VDD.n6644 VDD.n6643 0.731929
R5019 VDD.n6642 VDD.n6641 0.731929
R5020 VDD.n6640 VDD.n6639 0.731929
R5021 VDD.n6638 VDD.n6637 0.731929
R5022 VDD.n6636 VDD.n6635 0.731929
R5023 VDD.n6634 VDD.n6633 0.731929
R5024 VDD.n6632 VDD.n6631 0.731929
R5025 VDD.n6630 VDD.n6629 0.731929
R5026 VDD.n6628 VDD.n6627 0.731929
R5027 VDD.n6626 VDD.n6625 0.731929
R5028 VDD.n6624 VDD.n6623 0.731929
R5029 VDD.n6434 VDD.n6433 0.731929
R5030 VDD.n6436 VDD.n6435 0.731929
R5031 VDD.n6438 VDD.n6437 0.731929
R5032 VDD.n6440 VDD.n6439 0.731929
R5033 VDD.n6442 VDD.n6441 0.731929
R5034 VDD.n6444 VDD.n6443 0.731929
R5035 VDD.n6446 VDD.n6445 0.731929
R5036 VDD.n6448 VDD.n6447 0.731929
R5037 VDD.n6450 VDD.n6449 0.731929
R5038 VDD.n6452 VDD.n6451 0.731929
R5039 VDD.n6454 VDD.n6453 0.731929
R5040 VDD.n6456 VDD.n6455 0.731929
R5041 VDD.n6458 VDD.n6457 0.731929
R5042 VDD.n6460 VDD.n6459 0.731929
R5043 VDD.n6462 VDD.n6461 0.731929
R5044 VDD.n6464 VDD.n6463 0.731929
R5045 VDD.n6467 VDD.n6466 0.731929
R5046 VDD.n6471 VDD.n6469 0.731929
R5047 VDD.n6475 VDD.n6473 0.731929
R5048 VDD.n6479 VDD.n6477 0.731929
R5049 VDD.n6483 VDD.n6481 0.731929
R5050 VDD.n6390 VDD.n6389 0.72647
R5051 VDD.n6284 VDD.n6283 0.72647
R5052 VDD.n1794 VDD.n1374 0.718646
R5053 VDD.n805 VDD.n804 0.716028
R5054 VDD.n717 VDD.n716 0.716028
R5055 VDD.n629 VDD.n628 0.716028
R5056 VDD.n541 VDD.n540 0.716028
R5057 VDD.n453 VDD.n452 0.716028
R5058 VDD.n311 VDD.n310 0.698682
R5059 VDD.n6350 VDD.n6349 0.688261
R5060 VDD.n1616 VDD.n1612 0.65691
R5061 VDD.n1610 VDD.n1606 0.65691
R5062 VDD.n1604 VDD.n1600 0.65691
R5063 VDD.n1598 VDD.n1594 0.65691
R5064 VDD.n1592 VDD.n1588 0.65691
R5065 VDD.n1586 VDD.n1583 0.65691
R5066 VDD.n90 VDD.n89 0.647808
R5067 VDD.n3496 VDD.n3495 0.6405
R5068 VDD.n3540 VDD.n3539 0.6405
R5069 VDD.n3680 VDD.n3670 0.6405
R5070 VDD.n3848 VDD.n3847 0.6405
R5071 VDD.n3859 VDD.n3858 0.6405
R5072 VDD.n3899 VDD.n3898 0.6405
R5073 VDD.n3903 VDD.n3902 0.6405
R5074 VDD.n3997 VDD.n3996 0.6405
R5075 VDD.n4000 VDD.n3998 0.6405
R5076 VDD.n4023 VDD.n4021 0.6405
R5077 VDD.n4045 VDD.n4043 0.6405
R5078 VDD.n4064 VDD.n4062 0.6405
R5079 VDD.n4153 VDD.n4152 0.6405
R5080 VDD.n4194 VDD.n4193 0.6405
R5081 VDD.n4205 VDD.n4204 0.6405
R5082 VDD.n4220 VDD.n4219 0.6405
R5083 VDD.n4235 VDD.n4234 0.6405
R5084 VDD.n4239 VDD.n4238 0.6405
R5085 VDD.n4306 VDD.n4305 0.6405
R5086 VDD.n4327 VDD.n4326 0.6405
R5087 VDD.n4348 VDD.n4347 0.6405
R5088 VDD.n4367 VDD.n4366 0.6405
R5089 VDD.n4437 VDD.n4436 0.6405
R5090 VDD.n4477 VDD.n4476 0.6405
R5091 VDD.n4507 VDD.n4506 0.6405
R5092 VDD.n4546 VDD.n4545 0.6405
R5093 VDD.n4564 VDD.n4563 0.6405
R5094 VDD.n4567 VDD.n4566 0.6405
R5095 VDD.n4623 VDD.n4613 0.6405
R5096 VDD.n4786 VDD.n4785 0.6405
R5097 VDD.n4816 VDD.n4815 0.6405
R5098 VDD.n4834 VDD.n4822 0.6405
R5099 VDD.n4857 VDD.n4856 0.6405
R5100 VDD.n4884 VDD.n4883 0.6405
R5101 VDD.n4900 VDD.n4899 0.6405
R5102 VDD.n4923 VDD.n4922 0.6405
R5103 VDD.n5126 VDD.n5125 0.6405
R5104 VDD.n5268 VDD.n5267 0.6405
R5105 VDD.n1749 VDD.n1747 0.615885
R5106 VDD.n6396 VDD.n6395 0.573634
R5107 VDD.n6290 VDD.n6289 0.573634
R5108 VDD.n1208 VDD.n1207 0.56701
R5109 VDD.n785 VDD.n784 0.557022
R5110 VDD.n697 VDD.n696 0.557022
R5111 VDD.n609 VDD.n608 0.557022
R5112 VDD.n521 VDD.n520 0.557022
R5113 VDD.n433 VDD.n432 0.557022
R5114 VDD.n1189 VDD.n1104 0.554346
R5115 VDD.n1317 VDD.n1315 0.554346
R5116 VDD.n3010 VDD.t6 0.551225
R5117 VDD.n3014 VDD.n3013 0.551225
R5118 VDD.n3552 VDD.n3548 0.551225
R5119 VDD.n3678 VDD.n3677 0.551225
R5120 VDD.n3741 VDD.n3740 0.551225
R5121 VDD.n3913 VDD.n3909 0.551225
R5122 VDD.n4015 VDD.t72 0.551225
R5123 VDD.n4040 VDD.n4039 0.551225
R5124 VDD.n4094 VDD.n4093 0.551225
R5125 VDD.t135 VDD.n4111 0.551225
R5126 VDD.n4247 VDD.n4244 0.551225
R5127 VDD.n4362 VDD.n4361 0.551225
R5128 VDD.n4416 VDD.n4415 0.551225
R5129 VDD.t110 VDD.n4494 0.551225
R5130 VDD.n4579 VDD.n4575 0.551225
R5131 VDD.n4708 VDD.n4707 0.551225
R5132 VDD.n4766 VDD.n4765 0.551225
R5133 VDD.t2 VDD.n4805 0.551225
R5134 VDD.t83 VDD.n4895 0.551225
R5135 VDD.n4935 VDD.n4931 0.551225
R5136 VDD.n5062 VDD.n5061 0.551225
R5137 VDD.n5115 VDD.n5114 0.551225
R5138 VDD.n292 VDD.n291 0.54353
R5139 VDD.n6344 VDD.n6343 0.535425
R5140 VDD.n1206 VDD.n1205 0.533833
R5141 VDD.n1292 VDD.n1290 0.533833
R5142 VDD.n6696 VDD.n6621 0.528754
R5143 VDD.n6504 VDD.n6503 0.497216
R5144 VDD.n1755 VDD.n1751 0.492808
R5145 VDD.n1761 VDD.n1757 0.492808
R5146 VDD.n1767 VDD.n1763 0.492808
R5147 VDD.n1773 VDD.n1769 0.492808
R5148 VDD.n1779 VDD.n1775 0.492808
R5149 VDD.n1785 VDD.n1781 0.492808
R5150 VDD.n238 VDD.n237 0.465955
R5151 VDD.n253 VDD.n252 0.465955
R5152 VDD.n6697 VDD.n6696 0.455524
R5153 VDD.n1208 VDD.n114 0.455262
R5154 VDD.n900 VDD.n899 0.452265
R5155 VDD.n890 VDD.n889 0.452265
R5156 VDD.n1793 VDD.n1792 0.451782
R5157 VDD.n1581 VDD.n1579 0.451782
R5158 VDD.n1510 VDD.n1509 0.451782
R5159 VDD.n1524 VDD.n1523 0.431269
R5160 VDD.n3001 VDD.n2998 0.421259
R5161 VDD.n6402 VDD.n6401 0.420798
R5162 VDD.n6296 VDD.n6295 0.420798
R5163 VDD.n6713 VDD.n6710 0.420798
R5164 VDD.n1482 VDD.n1480 0.410756
R5165 VDD.n1487 VDD.n1485 0.410756
R5166 VDD.n1492 VDD.n1490 0.410756
R5167 VDD.n1497 VDD.n1495 0.410756
R5168 VDD.n1502 VDD.n1500 0.410756
R5169 VDD.n1507 VDD.n1505 0.410756
R5170 VDD.n2701 VDD.n2700 0.406849
R5171 VDD.n800 VDD.n799 0.398016
R5172 VDD.n712 VDD.n711 0.398016
R5173 VDD.n624 VDD.n623 0.398016
R5174 VDD.n536 VDD.n535 0.398016
R5175 VDD.n448 VDD.n447 0.398016
R5176 VDD.n306 VDD.n305 0.388379
R5177 VDD.n2651 VDD.n2647 0.383082
R5178 VDD.n2644 VDD.n2640 0.383082
R5179 VDD.n2637 VDD.n2633 0.383082
R5180 VDD.n2630 VDD.n2626 0.383082
R5181 VDD.n2623 VDD.n2619 0.383082
R5182 VDD.n2616 VDD.n2612 0.383082
R5183 VDD.n2609 VDD.n2605 0.383082
R5184 VDD.n2602 VDD.n2598 0.383082
R5185 VDD.n2595 VDD.n2591 0.383082
R5186 VDD.n2588 VDD.n2584 0.383082
R5187 VDD.n2581 VDD.n2577 0.383082
R5188 VDD.n2574 VDD.n2570 0.383082
R5189 VDD.n2567 VDD.n2563 0.383082
R5190 VDD.n2560 VDD.n2556 0.383082
R5191 VDD.n2553 VDD.n2549 0.383082
R5192 VDD.n2546 VDD.n2542 0.383082
R5193 VDD.n2539 VDD.n2535 0.383082
R5194 VDD.n2532 VDD.n2528 0.383082
R5195 VDD.n2525 VDD.n2521 0.383082
R5196 VDD.n2518 VDD.n2514 0.383082
R5197 VDD.n6338 VDD.n6337 0.38259
R5198 VDD.n2472 VDD.n2468 0.380364
R5199 VDD.n2465 VDD.n2461 0.380364
R5200 VDD.n2458 VDD.n2454 0.380364
R5201 VDD.n2451 VDD.n2447 0.380364
R5202 VDD.n2444 VDD.n2440 0.380364
R5203 VDD.n2437 VDD.n2433 0.380364
R5204 VDD.n2430 VDD.n2426 0.380364
R5205 VDD.n2423 VDD.n2419 0.380364
R5206 VDD.n2416 VDD.n2412 0.380364
R5207 VDD.n2409 VDD.n2405 0.380364
R5208 VDD.n2402 VDD.n2398 0.380364
R5209 VDD.n2395 VDD.n2391 0.380364
R5210 VDD.n2388 VDD.n2384 0.380364
R5211 VDD.n2381 VDD.n2377 0.380364
R5212 VDD.n2374 VDD.n2370 0.380364
R5213 VDD.n2367 VDD.n2363 0.380364
R5214 VDD.n2360 VDD.n2356 0.380364
R5215 VDD.n2353 VDD.n2349 0.380364
R5216 VDD.n2346 VDD.n2342 0.380364
R5217 VDD.n2339 VDD.n2335 0.380364
R5218 VDD.n94 VDD.n93 0.376971
R5219 VDD.n104 VDD.n103 0.376971
R5220 VDD.n875 VDD.n868 0.376971
R5221 VDD.n2293 VDD.n2289 0.375043
R5222 VDD.n2286 VDD.n2282 0.375043
R5223 VDD.n2279 VDD.n2275 0.375043
R5224 VDD.n2272 VDD.n2268 0.375043
R5225 VDD.n2265 VDD.n2261 0.375043
R5226 VDD.n2258 VDD.n2254 0.375043
R5227 VDD.n2251 VDD.n2247 0.375043
R5228 VDD.n2244 VDD.n2240 0.375043
R5229 VDD.n2237 VDD.n2233 0.375043
R5230 VDD.n2230 VDD.n2226 0.375043
R5231 VDD.n2223 VDD.n2219 0.375043
R5232 VDD.n2216 VDD.n2212 0.375043
R5233 VDD.n2209 VDD.n2205 0.375043
R5234 VDD.n2202 VDD.n2198 0.375043
R5235 VDD.n2195 VDD.n2191 0.375043
R5236 VDD.n2188 VDD.n2184 0.375043
R5237 VDD.n2181 VDD.n2177 0.375043
R5238 VDD.n2174 VDD.n2170 0.375043
R5239 VDD.n2167 VDD.n2163 0.375043
R5240 VDD.n2160 VDD.n2156 0.375043
R5241 VDD.n2114 VDD.n2113 0.373707
R5242 VDD.n2107 VDD.n2106 0.373707
R5243 VDD.n2100 VDD.n2099 0.373707
R5244 VDD.n2093 VDD.n2092 0.373707
R5245 VDD.n2086 VDD.n2085 0.373707
R5246 VDD.n2079 VDD.n2078 0.373707
R5247 VDD.n2072 VDD.n2071 0.373707
R5248 VDD.n2065 VDD.n2064 0.373707
R5249 VDD.n2058 VDD.n2057 0.373707
R5250 VDD.n2051 VDD.n2050 0.373707
R5251 VDD.n2044 VDD.n2043 0.373707
R5252 VDD.n2037 VDD.n2036 0.373707
R5253 VDD.n2030 VDD.n2029 0.373707
R5254 VDD.n2023 VDD.n2022 0.373707
R5255 VDD.n2016 VDD.n2015 0.373707
R5256 VDD.n2009 VDD.n2008 0.373707
R5257 VDD.n2002 VDD.n2001 0.373707
R5258 VDD.n1995 VDD.n1994 0.373707
R5259 VDD.n1988 VDD.n1987 0.373707
R5260 VDD.n1981 VDD.n1980 0.373707
R5261 VDD.n5854 VDD.n5853 0.369995
R5262 VDD.n5847 VDD.n5846 0.369995
R5263 VDD.n5840 VDD.n5839 0.369995
R5264 VDD.n5833 VDD.n5832 0.369995
R5265 VDD.n5826 VDD.n5825 0.369995
R5266 VDD.n5819 VDD.n5818 0.369995
R5267 VDD.n5812 VDD.n5811 0.369995
R5268 VDD.n5805 VDD.n5804 0.369995
R5269 VDD.n5798 VDD.n5797 0.369995
R5270 VDD.n5791 VDD.n5790 0.369995
R5271 VDD.n5784 VDD.n5783 0.369995
R5272 VDD.n5777 VDD.n5776 0.369995
R5273 VDD.n5770 VDD.n5769 0.369995
R5274 VDD.n5763 VDD.n5762 0.369995
R5275 VDD.n5756 VDD.n5755 0.369995
R5276 VDD.n5749 VDD.n5748 0.369995
R5277 VDD.n5742 VDD.n5741 0.369995
R5278 VDD.n5735 VDD.n5734 0.369995
R5279 VDD.n5728 VDD.n5727 0.369995
R5280 VDD.n5721 VDD.n5720 0.369995
R5281 VDD.n1935 VDD.n1934 0.369995
R5282 VDD.n1928 VDD.n1927 0.369995
R5283 VDD.n1921 VDD.n1920 0.369995
R5284 VDD.n1914 VDD.n1913 0.369995
R5285 VDD.n1907 VDD.n1906 0.369995
R5286 VDD.n1900 VDD.n1899 0.369995
R5287 VDD.n1893 VDD.n1892 0.369995
R5288 VDD.n1886 VDD.n1885 0.369995
R5289 VDD.n1879 VDD.n1878 0.369995
R5290 VDD.n1872 VDD.n1871 0.369995
R5291 VDD.n1865 VDD.n1864 0.369995
R5292 VDD.n1858 VDD.n1857 0.369995
R5293 VDD.n1851 VDD.n1850 0.369995
R5294 VDD.n1844 VDD.n1843 0.369995
R5295 VDD.n1837 VDD.n1836 0.369995
R5296 VDD.n1830 VDD.n1829 0.369995
R5297 VDD.n1823 VDD.n1822 0.369995
R5298 VDD.n1816 VDD.n1815 0.369995
R5299 VDD.n1809 VDD.n1808 0.369995
R5300 VDD.n1802 VDD.n1801 0.369995
R5301 VDD.n1621 VDD.n1620 0.369731
R5302 VDD.n5675 VDD.n5674 0.368684
R5303 VDD.n5668 VDD.n5667 0.368684
R5304 VDD.n5661 VDD.n5660 0.368684
R5305 VDD.n5654 VDD.n5653 0.368684
R5306 VDD.n5647 VDD.n5646 0.368684
R5307 VDD.n5640 VDD.n5639 0.368684
R5308 VDD.n5633 VDD.n5632 0.368684
R5309 VDD.n5626 VDD.n5625 0.368684
R5310 VDD.n5619 VDD.n5618 0.368684
R5311 VDD.n5612 VDD.n5611 0.368684
R5312 VDD.n5605 VDD.n5604 0.368684
R5313 VDD.n5598 VDD.n5597 0.368684
R5314 VDD.n5591 VDD.n5590 0.368684
R5315 VDD.n5584 VDD.n5583 0.368684
R5316 VDD.n5577 VDD.n5576 0.368684
R5317 VDD.n5570 VDD.n5569 0.368684
R5318 VDD.n5563 VDD.n5562 0.368684
R5319 VDD.n5556 VDD.n5555 0.368684
R5320 VDD.n5549 VDD.n5548 0.368684
R5321 VDD.n5542 VDD.n5541 0.368684
R5322 VDD.n3032 VDD.n3031 0.36765
R5323 VDD.n3503 VDD.n3501 0.36765
R5324 VDD.n3551 VDD.n3549 0.36765
R5325 VDD.n3701 VDD.t143 0.36765
R5326 VDD.n3719 VDD.n3718 0.36765
R5327 VDD.n3867 VDD.n3865 0.36765
R5328 VDD.n3912 VDD.n3910 0.36765
R5329 VDD.n3969 VDD.t11 0.36765
R5330 VDD.n4074 VDD.n4073 0.36765
R5331 VDD.n4209 VDD.n4208 0.36765
R5332 VDD.n4246 VDD.n4245 0.36765
R5333 VDD.n4395 VDD.n4394 0.36765
R5334 VDD.n4537 VDD.n4535 0.36765
R5335 VDD.n4578 VDD.n4576 0.36765
R5336 VDD.n4744 VDD.n4743 0.36765
R5337 VDD.n4891 VDD.n4889 0.36765
R5338 VDD.n5094 VDD.n5093 0.36765
R5339 VDD.n6033 VDD.n6032 0.360687
R5340 VDD.n6026 VDD.n6025 0.360687
R5341 VDD.n6019 VDD.n6018 0.360687
R5342 VDD.n6012 VDD.n6011 0.360687
R5343 VDD.n6005 VDD.n6004 0.360687
R5344 VDD.n5998 VDD.n5997 0.360687
R5345 VDD.n5991 VDD.n5990 0.360687
R5346 VDD.n5984 VDD.n5983 0.360687
R5347 VDD.n5977 VDD.n5976 0.360687
R5348 VDD.n5970 VDD.n5969 0.360687
R5349 VDD.n5963 VDD.n5962 0.360687
R5350 VDD.n5956 VDD.n5955 0.360687
R5351 VDD.n5949 VDD.n5948 0.360687
R5352 VDD.n5942 VDD.n5941 0.360687
R5353 VDD.n5935 VDD.n5934 0.360687
R5354 VDD.n5928 VDD.n5927 0.360687
R5355 VDD.n5921 VDD.n5920 0.360687
R5356 VDD.n5914 VDD.n5913 0.360687
R5357 VDD.n5907 VDD.n5906 0.360687
R5358 VDD.n5900 VDD.n5899 0.360687
R5359 VDD.n6212 VDD.n6211 0.35235
R5360 VDD.n6205 VDD.n6204 0.35235
R5361 VDD.n6198 VDD.n6197 0.35235
R5362 VDD.n6191 VDD.n6190 0.35235
R5363 VDD.n6184 VDD.n6183 0.35235
R5364 VDD.n6177 VDD.n6176 0.35235
R5365 VDD.n6170 VDD.n6169 0.35235
R5366 VDD.n6163 VDD.n6162 0.35235
R5367 VDD.n6156 VDD.n6155 0.35235
R5368 VDD.n6149 VDD.n6148 0.35235
R5369 VDD.n6142 VDD.n6141 0.35235
R5370 VDD.n6135 VDD.n6134 0.35235
R5371 VDD.n6128 VDD.n6127 0.35235
R5372 VDD.n6121 VDD.n6120 0.35235
R5373 VDD.n6114 VDD.n6113 0.35235
R5374 VDD.n6107 VDD.n6106 0.35235
R5375 VDD.n6100 VDD.n6099 0.35235
R5376 VDD.n6093 VDD.n6092 0.35235
R5377 VDD.n6086 VDD.n6085 0.35235
R5378 VDD.n6079 VDD.n6078 0.35235
R5379 VDD.n1312 VDD.n1309 0.349218
R5380 VDD.n1307 VDD.n1304 0.349218
R5381 VDD.n1302 VDD.n1299 0.349218
R5382 VDD.n1297 VDD.n1294 0.349218
R5383 VDD.n5496 VDD.n5495 0.346664
R5384 VDD.n5489 VDD.n5488 0.346664
R5385 VDD.n5482 VDD.n5481 0.346664
R5386 VDD.n5475 VDD.n5474 0.346664
R5387 VDD.n5468 VDD.n5467 0.346664
R5388 VDD.n5461 VDD.n5460 0.346664
R5389 VDD.n5454 VDD.n5453 0.346664
R5390 VDD.n5447 VDD.n5446 0.346664
R5391 VDD.n5440 VDD.n5439 0.346664
R5392 VDD.n5433 VDD.n5432 0.346664
R5393 VDD.n5426 VDD.n5425 0.346664
R5394 VDD.n5419 VDD.n5418 0.346664
R5395 VDD.n5412 VDD.n5411 0.346664
R5396 VDD.n5405 VDD.n5404 0.346664
R5397 VDD.n5398 VDD.n5397 0.346664
R5398 VDD.n5391 VDD.n5390 0.346664
R5399 VDD.n5384 VDD.n5383 0.346664
R5400 VDD.n5377 VDD.n5376 0.346664
R5401 VDD.n5370 VDD.n5369 0.346664
R5402 VDD.n5363 VDD.n5362 0.346664
R5403 VDD.n6430 VDD.n6429 0.344381
R5404 VDD.n1716 VDD.n1714 0.328705
R5405 VDD.n1721 VDD.n1719 0.328705
R5406 VDD.n1726 VDD.n1724 0.328705
R5407 VDD.n1732 VDD.n1730 0.328705
R5408 VDD.n1738 VDD.n1736 0.328705
R5409 VDD.n1744 VDD.n1742 0.328705
R5410 VDD.n1374 VDD.n1373 0.324592
R5411 VDD.n2997 VDD.n2834 0.3205
R5412 VDD.n3037 VDD.n3027 0.3205
R5413 VDD.n3516 VDD.n3515 0.3205
R5414 VDD.n3658 VDD.n3657 0.3205
R5415 VDD.n3690 VDD.n3688 0.3205
R5416 VDD.n3704 VDD.n3703 0.3205
R5417 VDD.n3724 VDD.n3714 0.3205
R5418 VDD.n4006 VDD.n4005 0.3205
R5419 VDD.n4029 VDD.n4028 0.3205
R5420 VDD.n4062 VDD.n4061 0.3205
R5421 VDD.n4078 VDD.n4070 0.3205
R5422 VDD.n4079 VDD.n4078 0.3205
R5423 VDD.n4158 VDD.n4157 0.3205
R5424 VDD.n4293 VDD.n4292 0.3205
R5425 VDD.n4311 VDD.n4310 0.3205
R5426 VDD.n4367 VDD.n4364 0.3205
R5427 VDD.n4383 VDD.n4382 0.3205
R5428 VDD.n4382 VDD.n4374 0.3205
R5429 VDD.n4399 VDD.n4391 0.3205
R5430 VDD.n4400 VDD.n4399 0.3205
R5431 VDD.n4460 VDD.n4459 0.3205
R5432 VDD.n4588 VDD.n4587 0.3205
R5433 VDD.n4608 VDD.n4607 0.3205
R5434 VDD.n4672 VDD.n4669 0.3205
R5435 VDD.n4692 VDD.n4691 0.3205
R5436 VDD.n4731 VDD.n4730 0.3205
R5437 VDD.n4730 VDD.n4720 0.3205
R5438 VDD.n4749 VDD.n4739 0.3205
R5439 VDD.n4750 VDD.n4749 0.3205
R5440 VDD.n4917 VDD.n4916 0.3205
R5441 VDD.n4983 VDD.n4980 0.3205
R5442 VDD.n4988 VDD.n4987 0.3205
R5443 VDD.n5005 VDD.n5004 0.3205
R5444 VDD.n5084 VDD.n5083 0.3205
R5445 VDD.n5083 VDD.n5075 0.3205
R5446 VDD.n5100 VDD.n5099 0.3205
R5447 VDD.n5099 VDD.n5098 0.3205
R5448 VDD.n5119 VDD.n5118 0.3205
R5449 VDD.n5140 VDD.n5139 0.3205
R5450 VDD.n5151 VDD.n5150 0.3205
R5451 VDD.n2704 VDD.n2703 0.29621
R5452 VDD.n2706 VDD.n2705 0.29621
R5453 VDD.n2708 VDD.n2707 0.29621
R5454 VDD.n2710 VDD.n2709 0.29621
R5455 VDD.n2712 VDD.n2711 0.29621
R5456 VDD.n2714 VDD.n2713 0.29621
R5457 VDD.n2716 VDD.n2715 0.29621
R5458 VDD.n2718 VDD.n2717 0.29621
R5459 VDD.n2720 VDD.n2719 0.29621
R5460 VDD.n2722 VDD.n2721 0.29621
R5461 VDD.n2724 VDD.n2723 0.29621
R5462 VDD.n2726 VDD.n2725 0.29621
R5463 VDD.n2728 VDD.n2727 0.29621
R5464 VDD.n2730 VDD.n2729 0.29621
R5465 VDD.n2733 VDD.n2731 0.29621
R5466 VDD.n2736 VDD.n2734 0.29621
R5467 VDD.n2739 VDD.n2737 0.29621
R5468 VDD.n2742 VDD.n2740 0.29621
R5469 VDD.n2745 VDD.n2743 0.29621
R5470 VDD.n2748 VDD.n2746 0.29621
R5471 VDD.n2751 VDD.n2749 0.29621
R5472 VDD.n2754 VDD.n2752 0.29621
R5473 VDD.n2757 VDD.n2755 0.29621
R5474 VDD.n2760 VDD.n2758 0.29621
R5475 VDD.n2763 VDD.n2761 0.29621
R5476 VDD.n2766 VDD.n2764 0.29621
R5477 VDD.n2769 VDD.n2767 0.29621
R5478 VDD.n2772 VDD.n2770 0.29621
R5479 VDD.n2775 VDD.n2773 0.29621
R5480 VDD.n2778 VDD.n2776 0.29621
R5481 VDD.n2781 VDD.n2779 0.29621
R5482 VDD.n2785 VDD.n2783 0.29621
R5483 VDD.n892 VDD.n158 0.279391
R5484 VDD.n1527 VDD.n1526 0.272099
R5485 VDD.n1529 VDD.n1528 0.270261
R5486 VDD.n6413 VDD.n6411 0.267963
R5487 VDD.n6407 VDD.n6405 0.267963
R5488 VDD.n6408 VDD.n6407 0.267963
R5489 VDD.n6401 VDD.n6399 0.267963
R5490 VDD.n6395 VDD.n6393 0.267963
R5491 VDD.n6389 VDD.n6387 0.267963
R5492 VDD.n6383 VDD.n6381 0.267963
R5493 VDD.n6375 VDD.n6373 0.267963
R5494 VDD.n6363 VDD.n6361 0.267963
R5495 VDD.n6355 VDD.n6353 0.267963
R5496 VDD.n6349 VDD.n6347 0.267963
R5497 VDD.n6343 VDD.n6341 0.267963
R5498 VDD.n6337 VDD.n6335 0.267963
R5499 VDD.n6331 VDD.n6329 0.267963
R5500 VDD.n6325 VDD.n6323 0.267963
R5501 VDD.n6307 VDD.n6305 0.267963
R5502 VDD.n6301 VDD.n6299 0.267963
R5503 VDD.n6302 VDD.n6301 0.267963
R5504 VDD.n6295 VDD.n6293 0.267963
R5505 VDD.n6289 VDD.n6287 0.267963
R5506 VDD.n6283 VDD.n6281 0.267963
R5507 VDD.n6277 VDD.n6275 0.267963
R5508 VDD.n6269 VDD.n6267 0.267963
R5509 VDD.n6258 VDD.n6256 0.267963
R5510 VDD.n5274 VDD.n5272 0.267963
R5511 VDD.n5278 VDD.n5276 0.267963
R5512 VDD.n1528 VDD.n1527 0.265665
R5513 VDD.n6709 VDD.n6708 0.253315
R5514 VDD.n6699 VDD.n6698 0.248811
R5515 VDD.n6700 VDD.n6699 0.248248
R5516 VDD.n1287 VDD.n1285 0.246654
R5517 VDD.n1282 VDD.n1280 0.246654
R5518 VDD.n1277 VDD.n1275 0.246654
R5519 VDD.n1272 VDD.n1270 0.246654
R5520 VDD.n1267 VDD.n1265 0.246654
R5521 VDD.n1262 VDD.n1260 0.246654
R5522 VDD.n6701 VDD.n6700 0.245432
R5523 VDD.n6705 VDD.n6704 0.245432
R5524 VDD.n6706 VDD.n6705 0.245432
R5525 VDD.n6707 VDD.n6706 0.245432
R5526 VDD.n6708 VDD.n6707 0.245432
R5527 VDD.n6702 VDD.n6701 0.239802
R5528 VDD.n876 VDD.n875 0.239009
R5529 VDD.n790 VDD.n789 0.239009
R5530 VDD.n702 VDD.n701 0.239009
R5531 VDD.n614 VDD.n613 0.239009
R5532 VDD.n526 VDD.n525 0.239009
R5533 VDD.n438 VDD.n437 0.239009
R5534 VDD.n6698 VDD.n6252 0.236869
R5535 VDD.n6699 VDD.n6073 0.236869
R5536 VDD.n6700 VDD.n5894 0.236869
R5537 VDD.n6701 VDD.n5715 0.236869
R5538 VDD.n6702 VDD.n5536 0.236869
R5539 VDD.n6704 VDD.n2691 0.236869
R5540 VDD.n6705 VDD.n2512 0.236869
R5541 VDD.n6706 VDD.n2333 0.236869
R5542 VDD.n6707 VDD.n2154 0.236869
R5543 VDD.n6708 VDD.n1975 0.236869
R5544 VDD.n6215 VDD.n6214 0.236284
R5545 VDD.n6217 VDD.n6216 0.236284
R5546 VDD.n6219 VDD.n6218 0.236284
R5547 VDD.n6221 VDD.n6220 0.236284
R5548 VDD.n6223 VDD.n6222 0.236284
R5549 VDD.n6225 VDD.n6224 0.236284
R5550 VDD.n6227 VDD.n6226 0.236284
R5551 VDD.n6229 VDD.n6228 0.236284
R5552 VDD.n6231 VDD.n6230 0.236284
R5553 VDD.n6233 VDD.n6232 0.236284
R5554 VDD.n6235 VDD.n6234 0.236284
R5555 VDD.n6237 VDD.n6236 0.236284
R5556 VDD.n6239 VDD.n6238 0.236284
R5557 VDD.n6241 VDD.n6240 0.236284
R5558 VDD.n6243 VDD.n6242 0.236284
R5559 VDD.n6245 VDD.n6244 0.236284
R5560 VDD.n6247 VDD.n6246 0.236284
R5561 VDD.n6249 VDD.n6248 0.236284
R5562 VDD.n6251 VDD.n6250 0.236284
R5563 VDD.n6036 VDD.n6035 0.236284
R5564 VDD.n6038 VDD.n6037 0.236284
R5565 VDD.n6040 VDD.n6039 0.236284
R5566 VDD.n6042 VDD.n6041 0.236284
R5567 VDD.n6044 VDD.n6043 0.236284
R5568 VDD.n6046 VDD.n6045 0.236284
R5569 VDD.n6048 VDD.n6047 0.236284
R5570 VDD.n6050 VDD.n6049 0.236284
R5571 VDD.n6052 VDD.n6051 0.236284
R5572 VDD.n6054 VDD.n6053 0.236284
R5573 VDD.n6056 VDD.n6055 0.236284
R5574 VDD.n6058 VDD.n6057 0.236284
R5575 VDD.n6060 VDD.n6059 0.236284
R5576 VDD.n6062 VDD.n6061 0.236284
R5577 VDD.n6064 VDD.n6063 0.236284
R5578 VDD.n6066 VDD.n6065 0.236284
R5579 VDD.n6068 VDD.n6067 0.236284
R5580 VDD.n6070 VDD.n6069 0.236284
R5581 VDD.n6072 VDD.n6071 0.236284
R5582 VDD.n5857 VDD.n5856 0.236284
R5583 VDD.n5859 VDD.n5858 0.236284
R5584 VDD.n5861 VDD.n5860 0.236284
R5585 VDD.n5863 VDD.n5862 0.236284
R5586 VDD.n5865 VDD.n5864 0.236284
R5587 VDD.n5867 VDD.n5866 0.236284
R5588 VDD.n5869 VDD.n5868 0.236284
R5589 VDD.n5871 VDD.n5870 0.236284
R5590 VDD.n5873 VDD.n5872 0.236284
R5591 VDD.n5875 VDD.n5874 0.236284
R5592 VDD.n5877 VDD.n5876 0.236284
R5593 VDD.n5879 VDD.n5878 0.236284
R5594 VDD.n5881 VDD.n5880 0.236284
R5595 VDD.n5883 VDD.n5882 0.236284
R5596 VDD.n5885 VDD.n5884 0.236284
R5597 VDD.n5887 VDD.n5886 0.236284
R5598 VDD.n5889 VDD.n5888 0.236284
R5599 VDD.n5891 VDD.n5890 0.236284
R5600 VDD.n5893 VDD.n5892 0.236284
R5601 VDD.n5678 VDD.n5677 0.236284
R5602 VDD.n5680 VDD.n5679 0.236284
R5603 VDD.n5682 VDD.n5681 0.236284
R5604 VDD.n5684 VDD.n5683 0.236284
R5605 VDD.n5686 VDD.n5685 0.236284
R5606 VDD.n5688 VDD.n5687 0.236284
R5607 VDD.n5690 VDD.n5689 0.236284
R5608 VDD.n5692 VDD.n5691 0.236284
R5609 VDD.n5694 VDD.n5693 0.236284
R5610 VDD.n5696 VDD.n5695 0.236284
R5611 VDD.n5698 VDD.n5697 0.236284
R5612 VDD.n5700 VDD.n5699 0.236284
R5613 VDD.n5702 VDD.n5701 0.236284
R5614 VDD.n5704 VDD.n5703 0.236284
R5615 VDD.n5706 VDD.n5705 0.236284
R5616 VDD.n5708 VDD.n5707 0.236284
R5617 VDD.n5710 VDD.n5709 0.236284
R5618 VDD.n5712 VDD.n5711 0.236284
R5619 VDD.n5714 VDD.n5713 0.236284
R5620 VDD.n5499 VDD.n5498 0.236284
R5621 VDD.n5501 VDD.n5500 0.236284
R5622 VDD.n5503 VDD.n5502 0.236284
R5623 VDD.n5505 VDD.n5504 0.236284
R5624 VDD.n5507 VDD.n5506 0.236284
R5625 VDD.n5509 VDD.n5508 0.236284
R5626 VDD.n5511 VDD.n5510 0.236284
R5627 VDD.n5513 VDD.n5512 0.236284
R5628 VDD.n5515 VDD.n5514 0.236284
R5629 VDD.n5517 VDD.n5516 0.236284
R5630 VDD.n5519 VDD.n5518 0.236284
R5631 VDD.n5521 VDD.n5520 0.236284
R5632 VDD.n5523 VDD.n5522 0.236284
R5633 VDD.n5525 VDD.n5524 0.236284
R5634 VDD.n5527 VDD.n5526 0.236284
R5635 VDD.n5529 VDD.n5528 0.236284
R5636 VDD.n5531 VDD.n5530 0.236284
R5637 VDD.n5533 VDD.n5532 0.236284
R5638 VDD.n5535 VDD.n5534 0.236284
R5639 VDD.n2654 VDD.n2653 0.236284
R5640 VDD.n2656 VDD.n2655 0.236284
R5641 VDD.n2658 VDD.n2657 0.236284
R5642 VDD.n2660 VDD.n2659 0.236284
R5643 VDD.n2662 VDD.n2661 0.236284
R5644 VDD.n2664 VDD.n2663 0.236284
R5645 VDD.n2666 VDD.n2665 0.236284
R5646 VDD.n2668 VDD.n2667 0.236284
R5647 VDD.n2670 VDD.n2669 0.236284
R5648 VDD.n2672 VDD.n2671 0.236284
R5649 VDD.n2674 VDD.n2673 0.236284
R5650 VDD.n2676 VDD.n2675 0.236284
R5651 VDD.n2678 VDD.n2677 0.236284
R5652 VDD.n2680 VDD.n2679 0.236284
R5653 VDD.n2682 VDD.n2681 0.236284
R5654 VDD.n2684 VDD.n2683 0.236284
R5655 VDD.n2686 VDD.n2685 0.236284
R5656 VDD.n2688 VDD.n2687 0.236284
R5657 VDD.n2690 VDD.n2689 0.236284
R5658 VDD.n2475 VDD.n2474 0.236284
R5659 VDD.n2477 VDD.n2476 0.236284
R5660 VDD.n2479 VDD.n2478 0.236284
R5661 VDD.n2481 VDD.n2480 0.236284
R5662 VDD.n2483 VDD.n2482 0.236284
R5663 VDD.n2485 VDD.n2484 0.236284
R5664 VDD.n2487 VDD.n2486 0.236284
R5665 VDD.n2489 VDD.n2488 0.236284
R5666 VDD.n2491 VDD.n2490 0.236284
R5667 VDD.n2493 VDD.n2492 0.236284
R5668 VDD.n2495 VDD.n2494 0.236284
R5669 VDD.n2497 VDD.n2496 0.236284
R5670 VDD.n2499 VDD.n2498 0.236284
R5671 VDD.n2501 VDD.n2500 0.236284
R5672 VDD.n2503 VDD.n2502 0.236284
R5673 VDD.n2505 VDD.n2504 0.236284
R5674 VDD.n2507 VDD.n2506 0.236284
R5675 VDD.n2509 VDD.n2508 0.236284
R5676 VDD.n2511 VDD.n2510 0.236284
R5677 VDD.n2296 VDD.n2295 0.236284
R5678 VDD.n2298 VDD.n2297 0.236284
R5679 VDD.n2300 VDD.n2299 0.236284
R5680 VDD.n2302 VDD.n2301 0.236284
R5681 VDD.n2304 VDD.n2303 0.236284
R5682 VDD.n2306 VDD.n2305 0.236284
R5683 VDD.n2308 VDD.n2307 0.236284
R5684 VDD.n2310 VDD.n2309 0.236284
R5685 VDD.n2312 VDD.n2311 0.236284
R5686 VDD.n2314 VDD.n2313 0.236284
R5687 VDD.n2316 VDD.n2315 0.236284
R5688 VDD.n2318 VDD.n2317 0.236284
R5689 VDD.n2320 VDD.n2319 0.236284
R5690 VDD.n2322 VDD.n2321 0.236284
R5691 VDD.n2324 VDD.n2323 0.236284
R5692 VDD.n2326 VDD.n2325 0.236284
R5693 VDD.n2328 VDD.n2327 0.236284
R5694 VDD.n2330 VDD.n2329 0.236284
R5695 VDD.n2332 VDD.n2331 0.236284
R5696 VDD.n2117 VDD.n2116 0.236284
R5697 VDD.n2119 VDD.n2118 0.236284
R5698 VDD.n2121 VDD.n2120 0.236284
R5699 VDD.n2123 VDD.n2122 0.236284
R5700 VDD.n2125 VDD.n2124 0.236284
R5701 VDD.n2127 VDD.n2126 0.236284
R5702 VDD.n2129 VDD.n2128 0.236284
R5703 VDD.n2131 VDD.n2130 0.236284
R5704 VDD.n2133 VDD.n2132 0.236284
R5705 VDD.n2135 VDD.n2134 0.236284
R5706 VDD.n2137 VDD.n2136 0.236284
R5707 VDD.n2139 VDD.n2138 0.236284
R5708 VDD.n2141 VDD.n2140 0.236284
R5709 VDD.n2143 VDD.n2142 0.236284
R5710 VDD.n2145 VDD.n2144 0.236284
R5711 VDD.n2147 VDD.n2146 0.236284
R5712 VDD.n2149 VDD.n2148 0.236284
R5713 VDD.n2151 VDD.n2150 0.236284
R5714 VDD.n2153 VDD.n2152 0.236284
R5715 VDD.n1938 VDD.n1937 0.236284
R5716 VDD.n1940 VDD.n1939 0.236284
R5717 VDD.n1942 VDD.n1941 0.236284
R5718 VDD.n1944 VDD.n1943 0.236284
R5719 VDD.n1946 VDD.n1945 0.236284
R5720 VDD.n1948 VDD.n1947 0.236284
R5721 VDD.n1950 VDD.n1949 0.236284
R5722 VDD.n1952 VDD.n1951 0.236284
R5723 VDD.n1954 VDD.n1953 0.236284
R5724 VDD.n1956 VDD.n1955 0.236284
R5725 VDD.n1958 VDD.n1957 0.236284
R5726 VDD.n1960 VDD.n1959 0.236284
R5727 VDD.n1962 VDD.n1961 0.236284
R5728 VDD.n1964 VDD.n1963 0.236284
R5729 VDD.n1966 VDD.n1965 0.236284
R5730 VDD.n1968 VDD.n1967 0.236284
R5731 VDD.n1970 VDD.n1969 0.236284
R5732 VDD.n1972 VDD.n1971 0.236284
R5733 VDD.n1974 VDD.n1973 0.236284
R5734 VDD.n1373 VDD.n1372 0.236249
R5735 VDD.n296 VDD.n295 0.233227
R5736 VDD.n6704 VDD.n6703 0.231919
R5737 VDD.n6420 VDD.n6417 0.229754
R5738 VDD.n6332 VDD.n6331 0.229754
R5739 VDD.n6314 VDD.n6311 0.229754
R5740 VDD.n1525 VDD.n1524 0.21053
R5741 VDD.n1790 VDD.n1789 0.205628
R5742 VDD.n6696 VDD.n6695 0.203675
R5743 VDD.n6498 VDD.n6497 0.191545
R5744 VDD.n6426 VDD.n6425 0.191545
R5745 VDD.n6320 VDD.n6319 0.191545
R5746 VDD.n2995 VDD.n2994 0.184075
R5747 VDD.n3035 VDD.n3034 0.184075
R5748 VDD.t61 VDD.n3418 0.184075
R5749 VDD.t88 VDD.n3551 0.184075
R5750 VDD.n3701 VDD.n3700 0.184075
R5751 VDD.n3722 VDD.n3721 0.184075
R5752 VDD.n3842 VDD.t0 0.184075
R5753 VDD.n4059 VDD.n4058 0.184075
R5754 VDD.n4076 VDD.n4075 0.184075
R5755 VDD.n4380 VDD.n4379 0.184075
R5756 VDD.n4397 VDD.n4396 0.184075
R5757 VDD.t115 VDD.n4617 0.184075
R5758 VDD.n4728 VDD.n4727 0.184075
R5759 VDD.n4747 VDD.n4746 0.184075
R5760 VDD.n4762 VDD.t8 0.184075
R5761 VDD.n4934 VDD.t98 0.184075
R5762 VDD.t98 VDD.n4932 0.184075
R5763 VDD.t120 VDD.n5081 0.184075
R5764 VDD.n5096 VDD.n5095 0.184075
R5765 VDD.n1576 VDD.n1574 0.164603
R5766 VDD.n1450 VDD.n1447 0.164603
R5767 VDD.n1455 VDD.n1452 0.164603
R5768 VDD.n1460 VDD.n1457 0.164603
R5769 VDD.n1465 VDD.n1462 0.164603
R5770 VDD.n1470 VDD.n1467 0.164603
R5771 VDD.n879 VDD.n878 0.158109
R5772 VDD.n243 VDD.n242 0.155652
R5773 VDD.n248 VDD.n247 0.155652
R5774 VDD.n132 VDD.n131 0.151088
R5775 VDD.n120 VDD.n119 0.151088
R5776 VDD.n1320 VDD.n1221 0.14409
R5777 VDD.n1524 VDD.n1515 0.14409
R5778 VDD.n1526 VDD.n1525 0.131714
R5779 VDD.n1372 VDD.n1320 0.125175
R5780 VDD.n1475 VDD.n1473 0.123577
R5781 VDD VDD.n6791 0.120996
R5782 VDD.n6703 VDD.n6702 0.11818
R5783 VDD.n6414 VDD.n6413 0.115127
R5784 VDD.n6308 VDD.n6307 0.115127
R5785 VDD.n6703 VDD.n5357 0.0984167
R5786 VDD.n1661 VDD.n1529 0.094394
R5787 VDD.n6709 VDD.n1796 0.0916052
R5788 VDD.n3051 VDD.n3050 0.088
R5789 VDD.n3054 VDD.n3053 0.088
R5790 VDD.n3068 VDD.n3067 0.088
R5791 VDD.n3082 VDD.n3081 0.088
R5792 VDD.n3085 VDD.n3084 0.088
R5793 VDD.n3099 VDD.n3098 0.088
R5794 VDD.n3113 VDD.n3112 0.088
R5795 VDD.n3116 VDD.n3115 0.088
R5796 VDD.n3130 VDD.n3129 0.088
R5797 VDD.n3144 VDD.n3143 0.088
R5798 VDD.n3147 VDD.n3146 0.088
R5799 VDD.n3161 VDD.n3160 0.088
R5800 VDD.n3175 VDD.n3174 0.088
R5801 VDD.n3178 VDD.n3177 0.088
R5802 VDD.n3192 VDD.n3191 0.088
R5803 VDD.n3206 VDD.n3205 0.088
R5804 VDD.n3209 VDD.n3208 0.088
R5805 VDD.n3223 VDD.n3222 0.088
R5806 VDD.n3237 VDD.n3236 0.088
R5807 VDD.n3240 VDD.n3239 0.088
R5808 VDD.n3254 VDD.n3253 0.088
R5809 VDD.n3268 VDD.n3267 0.088
R5810 VDD.n3271 VDD.n3270 0.088
R5811 VDD.n3285 VDD.n3284 0.088
R5812 VDD.n3299 VDD.n3298 0.088
R5813 VDD.n3302 VDD.n3301 0.088
R5814 VDD.n3316 VDD.n3315 0.088
R5815 VDD.n3330 VDD.n3329 0.088
R5816 VDD.n3333 VDD.n3332 0.088
R5817 VDD.n3347 VDD.n3346 0.088
R5818 VDD.n3361 VDD.n3360 0.088
R5819 VDD.n3364 VDD.n3363 0.088
R5820 VDD.n3378 VDD.n3377 0.088
R5821 VDD.n4229 VDD.n4223 0.088
R5822 VDD.n4068 VDD.n4067 0.0859167
R5823 VDD.n367 VDD.n361 0.0856449
R5824 VDD.n3897 VDD.n3896 0.0838333
R5825 VDD.n1659 VDD.n1655 0.0825513
R5826 VDD.n1653 VDD.n1649 0.0825513
R5827 VDD.n1647 VDD.n1643 0.0825513
R5828 VDD.n1641 VDD.n1637 0.0825513
R5829 VDD.n1635 VDD.n1631 0.0825513
R5830 VDD.n1629 VDD.n1625 0.0825513
R5831 VDD.n3731 VDD.n3730 0.08175
R5832 VDD.n795 VDD.n794 0.0800031
R5833 VDD.n707 VDD.n706 0.0800031
R5834 VDD.n619 VDD.n618 0.0800031
R5835 VDD.n531 VDD.n530 0.0800031
R5836 VDD.n443 VDD.n442 0.0800031
R5837 VDD.n3560 VDD.n3559 0.0796667
R5838 VDD.n301 VDD.n300 0.0780758
R5839 VDD.n3003 VDD.n3002 0.0775833
R5840 VDD.n6426 VDD.n6423 0.0769179
R5841 VDD.n6326 VDD.n6325 0.0769179
R5842 VDD.n6320 VDD.n6317 0.0769179
R5843 VDD.n6505 VDD.n6431 0.0692023
R5844 VDD.n6431 VDD.n6427 0.0692023
R5845 VDD.n6427 VDD.n6421 0.0692023
R5846 VDD.n6421 VDD.n6415 0.0692023
R5847 VDD.n6415 VDD.n6409 0.0692023
R5848 VDD.n6409 VDD.n6403 0.0692023
R5849 VDD.n6403 VDD.n6397 0.0692023
R5850 VDD.n6397 VDD.n6391 0.0692023
R5851 VDD.n6391 VDD.n6385 0.0692023
R5852 VDD.n6385 VDD.n6379 0.0692023
R5853 VDD.n6379 VDD.n6371 0.0692023
R5854 VDD.n6371 VDD.n6365 0.0692023
R5855 VDD.n6365 VDD.n6357 0.0692023
R5856 VDD.n6357 VDD.n6351 0.0692023
R5857 VDD.n6351 VDD.n6345 0.0692023
R5858 VDD.n6345 VDD.n6339 0.0692023
R5859 VDD.n6339 VDD.n6333 0.0692023
R5860 VDD.n6333 VDD.n6327 0.0692023
R5861 VDD.n6327 VDD.n6321 0.0692023
R5862 VDD.n6321 VDD.n6315 0.0692023
R5863 VDD.n6315 VDD.n6309 0.0692023
R5864 VDD.n6309 VDD.n6303 0.0692023
R5865 VDD.n6303 VDD.n6297 0.0692023
R5866 VDD.n6297 VDD.n6291 0.0692023
R5867 VDD.n6291 VDD.n6285 0.0692023
R5868 VDD.n6285 VDD.n6279 0.0692023
R5869 VDD.n6279 VDD.n6273 0.0692023
R5870 VDD.n6273 VDD.n6265 0.0692023
R5871 VDD.n186 VDD.n181 0.0657174
R5872 VDD.n191 VDD.n186 0.0657174
R5873 VDD.n196 VDD.n191 0.0657174
R5874 VDD.n204 VDD.n196 0.0657174
R5875 VDD.n209 VDD.n204 0.0657174
R5876 VDD.n214 VDD.n209 0.0657174
R5877 VDD.n219 VDD.n214 0.0657174
R5878 VDD.n224 VDD.n219 0.0657174
R5879 VDD.n229 VDD.n224 0.0657174
R5880 VDD.n234 VDD.n229 0.0657174
R5881 VDD.n239 VDD.n234 0.0657174
R5882 VDD.n244 VDD.n239 0.0657174
R5883 VDD.n249 VDD.n244 0.0657174
R5884 VDD.n254 VDD.n249 0.0657174
R5885 VDD.n259 VDD.n254 0.0657174
R5886 VDD.n260 VDD.n259 0.0657174
R5887 VDD.n302 VDD.n297 0.0657174
R5888 VDD.n307 VDD.n302 0.0657174
R5889 VDD.n312 VDD.n307 0.0657174
R5890 VDD.n317 VDD.n312 0.0657174
R5891 VDD.n322 VDD.n317 0.0657174
R5892 VDD.n327 VDD.n322 0.0657174
R5893 VDD.n332 VDD.n327 0.0657174
R5894 VDD.n337 VDD.n332 0.0657174
R5895 VDD.n345 VDD.n337 0.0657174
R5896 VDD.n350 VDD.n345 0.0657174
R5897 VDD.n355 VDD.n350 0.0657174
R5898 VDD.n361 VDD.n355 0.0657174
R5899 VDD.n878 VDD.n877 0.0657174
R5900 VDD.n877 VDD.n864 0.0657174
R5901 VDD.n864 VDD.n859 0.0657174
R5902 VDD.n859 VDD.n854 0.0657174
R5903 VDD.n854 VDD.n849 0.0657174
R5904 VDD.n849 VDD.n844 0.0657174
R5905 VDD.n844 VDD.n839 0.0657174
R5906 VDD.n839 VDD.n831 0.0657174
R5907 VDD.n831 VDD.n826 0.0657174
R5908 VDD.n826 VDD.n821 0.0657174
R5909 VDD.n821 VDD.n816 0.0657174
R5910 VDD.n816 VDD.n811 0.0657174
R5911 VDD.n811 VDD.n806 0.0657174
R5912 VDD.n806 VDD.n801 0.0657174
R5913 VDD.n801 VDD.n796 0.0657174
R5914 VDD.n796 VDD.n791 0.0657174
R5915 VDD.n791 VDD.n786 0.0657174
R5916 VDD.n786 VDD.n781 0.0657174
R5917 VDD.n781 VDD.n776 0.0657174
R5918 VDD.n776 VDD.n771 0.0657174
R5919 VDD.n771 VDD.n766 0.0657174
R5920 VDD.n766 VDD.n761 0.0657174
R5921 VDD.n761 VDD.n756 0.0657174
R5922 VDD.n756 VDD.n751 0.0657174
R5923 VDD.n751 VDD.n743 0.0657174
R5924 VDD.n743 VDD.n738 0.0657174
R5925 VDD.n738 VDD.n733 0.0657174
R5926 VDD.n733 VDD.n728 0.0657174
R5927 VDD.n728 VDD.n723 0.0657174
R5928 VDD.n723 VDD.n718 0.0657174
R5929 VDD.n718 VDD.n713 0.0657174
R5930 VDD.n713 VDD.n708 0.0657174
R5931 VDD.n708 VDD.n703 0.0657174
R5932 VDD.n703 VDD.n698 0.0657174
R5933 VDD.n698 VDD.n693 0.0657174
R5934 VDD.n693 VDD.n688 0.0657174
R5935 VDD.n688 VDD.n683 0.0657174
R5936 VDD.n683 VDD.n678 0.0657174
R5937 VDD.n678 VDD.n673 0.0657174
R5938 VDD.n673 VDD.n668 0.0657174
R5939 VDD.n668 VDD.n663 0.0657174
R5940 VDD.n663 VDD.n655 0.0657174
R5941 VDD.n655 VDD.n650 0.0657174
R5942 VDD.n650 VDD.n645 0.0657174
R5943 VDD.n645 VDD.n640 0.0657174
R5944 VDD.n640 VDD.n635 0.0657174
R5945 VDD.n635 VDD.n630 0.0657174
R5946 VDD.n630 VDD.n625 0.0657174
R5947 VDD.n625 VDD.n620 0.0657174
R5948 VDD.n620 VDD.n615 0.0657174
R5949 VDD.n615 VDD.n610 0.0657174
R5950 VDD.n610 VDD.n605 0.0657174
R5951 VDD.n605 VDD.n600 0.0657174
R5952 VDD.n600 VDD.n595 0.0657174
R5953 VDD.n595 VDD.n590 0.0657174
R5954 VDD.n590 VDD.n585 0.0657174
R5955 VDD.n585 VDD.n580 0.0657174
R5956 VDD.n580 VDD.n575 0.0657174
R5957 VDD.n575 VDD.n567 0.0657174
R5958 VDD.n567 VDD.n562 0.0657174
R5959 VDD.n562 VDD.n557 0.0657174
R5960 VDD.n557 VDD.n552 0.0657174
R5961 VDD.n552 VDD.n547 0.0657174
R5962 VDD.n547 VDD.n542 0.0657174
R5963 VDD.n542 VDD.n537 0.0657174
R5964 VDD.n537 VDD.n532 0.0657174
R5965 VDD.n532 VDD.n527 0.0657174
R5966 VDD.n527 VDD.n522 0.0657174
R5967 VDD.n522 VDD.n517 0.0657174
R5968 VDD.n517 VDD.n512 0.0657174
R5969 VDD.n512 VDD.n507 0.0657174
R5970 VDD.n507 VDD.n502 0.0657174
R5971 VDD.n502 VDD.n497 0.0657174
R5972 VDD.n497 VDD.n492 0.0657174
R5973 VDD.n492 VDD.n487 0.0657174
R5974 VDD.n487 VDD.n479 0.0657174
R5975 VDD.n479 VDD.n474 0.0657174
R5976 VDD.n474 VDD.n469 0.0657174
R5977 VDD.n469 VDD.n464 0.0657174
R5978 VDD.n464 VDD.n459 0.0657174
R5979 VDD.n459 VDD.n454 0.0657174
R5980 VDD.n454 VDD.n449 0.0657174
R5981 VDD.n449 VDD.n444 0.0657174
R5982 VDD.n444 VDD.n439 0.0657174
R5983 VDD.n439 VDD.n434 0.0657174
R5984 VDD.n434 VDD.n429 0.0657174
R5985 VDD.n429 VDD.n424 0.0657174
R5986 VDD.n424 VDD.n419 0.0657174
R5987 VDD.n419 VDD.n414 0.0657174
R5988 VDD.n414 VDD.n409 0.0657174
R5989 VDD.n409 VDD.n404 0.0657174
R5990 VDD.n404 VDD.n399 0.0657174
R5991 VDD.n399 VDD.n391 0.0657174
R5992 VDD.n391 VDD.n386 0.0657174
R5993 VDD.n386 VDD.n381 0.0657174
R5994 VDD.n381 VDD.n376 0.0657174
R5995 VDD.n376 VDD.n367 0.0657174
R5996 VDD.n1018 VDD.n947 0.0657174
R5997 VDD.n947 VDD.n942 0.0657174
R5998 VDD.n942 VDD.n937 0.0657174
R5999 VDD.n937 VDD.n932 0.0657174
R6000 VDD.n932 VDD.n927 0.0657174
R6001 VDD.n927 VDD.n922 0.0657174
R6002 VDD.n922 VDD.n914 0.0657174
R6003 VDD.n914 VDD.n909 0.0657174
R6004 VDD.n909 VDD.n904 0.0657174
R6005 VDD.n5031 VDD.n5030 0.063
R6006 VDD.n904 VDD.n902 0.0620942
R6007 VDD.n4862 VDD.n4861 0.0609167
R6008 VDD.n4697 VDD.n4696 0.0588333
R6009 VDD.n4531 VDD.n4530 0.05675
R6010 VDD.n4372 VDD.n4370 0.0546667
R6011 VDD.n6216 VDD.n6215 0.0527417
R6012 VDD.n6218 VDD.n6217 0.0527417
R6013 VDD.n6220 VDD.n6219 0.0527417
R6014 VDD.n6222 VDD.n6221 0.0527417
R6015 VDD.n6224 VDD.n6223 0.0527417
R6016 VDD.n6226 VDD.n6225 0.0527417
R6017 VDD.n6228 VDD.n6227 0.0527417
R6018 VDD.n6230 VDD.n6229 0.0527417
R6019 VDD.n6232 VDD.n6231 0.0527417
R6020 VDD.n6234 VDD.n6233 0.0527417
R6021 VDD.n6236 VDD.n6235 0.0527417
R6022 VDD.n6238 VDD.n6237 0.0527417
R6023 VDD.n6240 VDD.n6239 0.0527417
R6024 VDD.n6242 VDD.n6241 0.0527417
R6025 VDD.n6244 VDD.n6243 0.0527417
R6026 VDD.n6246 VDD.n6245 0.0527417
R6027 VDD.n6248 VDD.n6247 0.0527417
R6028 VDD.n6250 VDD.n6249 0.0527417
R6029 VDD.n6252 VDD.n6251 0.0527417
R6030 VDD.n6037 VDD.n6036 0.0527417
R6031 VDD.n6039 VDD.n6038 0.0527417
R6032 VDD.n6041 VDD.n6040 0.0527417
R6033 VDD.n6043 VDD.n6042 0.0527417
R6034 VDD.n6045 VDD.n6044 0.0527417
R6035 VDD.n6047 VDD.n6046 0.0527417
R6036 VDD.n6049 VDD.n6048 0.0527417
R6037 VDD.n6051 VDD.n6050 0.0527417
R6038 VDD.n6053 VDD.n6052 0.0527417
R6039 VDD.n6055 VDD.n6054 0.0527417
R6040 VDD.n6057 VDD.n6056 0.0527417
R6041 VDD.n6059 VDD.n6058 0.0527417
R6042 VDD.n6061 VDD.n6060 0.0527417
R6043 VDD.n6063 VDD.n6062 0.0527417
R6044 VDD.n6065 VDD.n6064 0.0527417
R6045 VDD.n6067 VDD.n6066 0.0527417
R6046 VDD.n6069 VDD.n6068 0.0527417
R6047 VDD.n6071 VDD.n6070 0.0527417
R6048 VDD.n6073 VDD.n6072 0.0527417
R6049 VDD.n5858 VDD.n5857 0.0527417
R6050 VDD.n5860 VDD.n5859 0.0527417
R6051 VDD.n5862 VDD.n5861 0.0527417
R6052 VDD.n5864 VDD.n5863 0.0527417
R6053 VDD.n5866 VDD.n5865 0.0527417
R6054 VDD.n5868 VDD.n5867 0.0527417
R6055 VDD.n5870 VDD.n5869 0.0527417
R6056 VDD.n5872 VDD.n5871 0.0527417
R6057 VDD.n5874 VDD.n5873 0.0527417
R6058 VDD.n5876 VDD.n5875 0.0527417
R6059 VDD.n5878 VDD.n5877 0.0527417
R6060 VDD.n5880 VDD.n5879 0.0527417
R6061 VDD.n5882 VDD.n5881 0.0527417
R6062 VDD.n5884 VDD.n5883 0.0527417
R6063 VDD.n5886 VDD.n5885 0.0527417
R6064 VDD.n5888 VDD.n5887 0.0527417
R6065 VDD.n5890 VDD.n5889 0.0527417
R6066 VDD.n5892 VDD.n5891 0.0527417
R6067 VDD.n5894 VDD.n5893 0.0527417
R6068 VDD.n5679 VDD.n5678 0.0527417
R6069 VDD.n5681 VDD.n5680 0.0527417
R6070 VDD.n5683 VDD.n5682 0.0527417
R6071 VDD.n5685 VDD.n5684 0.0527417
R6072 VDD.n5687 VDD.n5686 0.0527417
R6073 VDD.n5689 VDD.n5688 0.0527417
R6074 VDD.n5691 VDD.n5690 0.0527417
R6075 VDD.n5693 VDD.n5692 0.0527417
R6076 VDD.n5695 VDD.n5694 0.0527417
R6077 VDD.n5697 VDD.n5696 0.0527417
R6078 VDD.n5699 VDD.n5698 0.0527417
R6079 VDD.n5701 VDD.n5700 0.0527417
R6080 VDD.n5703 VDD.n5702 0.0527417
R6081 VDD.n5705 VDD.n5704 0.0527417
R6082 VDD.n5707 VDD.n5706 0.0527417
R6083 VDD.n5709 VDD.n5708 0.0527417
R6084 VDD.n5711 VDD.n5710 0.0527417
R6085 VDD.n5713 VDD.n5712 0.0527417
R6086 VDD.n5715 VDD.n5714 0.0527417
R6087 VDD.n5500 VDD.n5499 0.0527417
R6088 VDD.n5502 VDD.n5501 0.0527417
R6089 VDD.n5504 VDD.n5503 0.0527417
R6090 VDD.n5506 VDD.n5505 0.0527417
R6091 VDD.n5508 VDD.n5507 0.0527417
R6092 VDD.n5510 VDD.n5509 0.0527417
R6093 VDD.n5512 VDD.n5511 0.0527417
R6094 VDD.n5514 VDD.n5513 0.0527417
R6095 VDD.n5516 VDD.n5515 0.0527417
R6096 VDD.n5518 VDD.n5517 0.0527417
R6097 VDD.n5520 VDD.n5519 0.0527417
R6098 VDD.n5522 VDD.n5521 0.0527417
R6099 VDD.n5524 VDD.n5523 0.0527417
R6100 VDD.n5526 VDD.n5525 0.0527417
R6101 VDD.n5528 VDD.n5527 0.0527417
R6102 VDD.n5530 VDD.n5529 0.0527417
R6103 VDD.n5532 VDD.n5531 0.0527417
R6104 VDD.n5534 VDD.n5533 0.0527417
R6105 VDD.n5536 VDD.n5535 0.0527417
R6106 VDD.n2655 VDD.n2654 0.0527417
R6107 VDD.n2657 VDD.n2656 0.0527417
R6108 VDD.n2659 VDD.n2658 0.0527417
R6109 VDD.n2661 VDD.n2660 0.0527417
R6110 VDD.n2663 VDD.n2662 0.0527417
R6111 VDD.n2665 VDD.n2664 0.0527417
R6112 VDD.n2667 VDD.n2666 0.0527417
R6113 VDD.n2669 VDD.n2668 0.0527417
R6114 VDD.n2671 VDD.n2670 0.0527417
R6115 VDD.n2673 VDD.n2672 0.0527417
R6116 VDD.n2675 VDD.n2674 0.0527417
R6117 VDD.n2677 VDD.n2676 0.0527417
R6118 VDD.n2679 VDD.n2678 0.0527417
R6119 VDD.n2681 VDD.n2680 0.0527417
R6120 VDD.n2683 VDD.n2682 0.0527417
R6121 VDD.n2685 VDD.n2684 0.0527417
R6122 VDD.n2687 VDD.n2686 0.0527417
R6123 VDD.n2689 VDD.n2688 0.0527417
R6124 VDD.n2691 VDD.n2690 0.0527417
R6125 VDD.n2476 VDD.n2475 0.0527417
R6126 VDD.n2478 VDD.n2477 0.0527417
R6127 VDD.n2480 VDD.n2479 0.0527417
R6128 VDD.n2482 VDD.n2481 0.0527417
R6129 VDD.n2484 VDD.n2483 0.0527417
R6130 VDD.n2486 VDD.n2485 0.0527417
R6131 VDD.n2488 VDD.n2487 0.0527417
R6132 VDD.n2490 VDD.n2489 0.0527417
R6133 VDD.n2492 VDD.n2491 0.0527417
R6134 VDD.n2494 VDD.n2493 0.0527417
R6135 VDD.n2496 VDD.n2495 0.0527417
R6136 VDD.n2498 VDD.n2497 0.0527417
R6137 VDD.n2500 VDD.n2499 0.0527417
R6138 VDD.n2502 VDD.n2501 0.0527417
R6139 VDD.n2504 VDD.n2503 0.0527417
R6140 VDD.n2506 VDD.n2505 0.0527417
R6141 VDD.n2508 VDD.n2507 0.0527417
R6142 VDD.n2510 VDD.n2509 0.0527417
R6143 VDD.n2512 VDD.n2511 0.0527417
R6144 VDD.n2297 VDD.n2296 0.0527417
R6145 VDD.n2299 VDD.n2298 0.0527417
R6146 VDD.n2301 VDD.n2300 0.0527417
R6147 VDD.n2303 VDD.n2302 0.0527417
R6148 VDD.n2305 VDD.n2304 0.0527417
R6149 VDD.n2307 VDD.n2306 0.0527417
R6150 VDD.n2309 VDD.n2308 0.0527417
R6151 VDD.n2311 VDD.n2310 0.0527417
R6152 VDD.n2313 VDD.n2312 0.0527417
R6153 VDD.n2315 VDD.n2314 0.0527417
R6154 VDD.n2317 VDD.n2316 0.0527417
R6155 VDD.n2319 VDD.n2318 0.0527417
R6156 VDD.n2321 VDD.n2320 0.0527417
R6157 VDD.n2323 VDD.n2322 0.0527417
R6158 VDD.n2325 VDD.n2324 0.0527417
R6159 VDD.n2327 VDD.n2326 0.0527417
R6160 VDD.n2329 VDD.n2328 0.0527417
R6161 VDD.n2331 VDD.n2330 0.0527417
R6162 VDD.n2333 VDD.n2332 0.0527417
R6163 VDD.n2118 VDD.n2117 0.0527417
R6164 VDD.n2120 VDD.n2119 0.0527417
R6165 VDD.n2122 VDD.n2121 0.0527417
R6166 VDD.n2124 VDD.n2123 0.0527417
R6167 VDD.n2126 VDD.n2125 0.0527417
R6168 VDD.n2128 VDD.n2127 0.0527417
R6169 VDD.n2130 VDD.n2129 0.0527417
R6170 VDD.n2132 VDD.n2131 0.0527417
R6171 VDD.n2134 VDD.n2133 0.0527417
R6172 VDD.n2136 VDD.n2135 0.0527417
R6173 VDD.n2138 VDD.n2137 0.0527417
R6174 VDD.n2140 VDD.n2139 0.0527417
R6175 VDD.n2142 VDD.n2141 0.0527417
R6176 VDD.n2144 VDD.n2143 0.0527417
R6177 VDD.n2146 VDD.n2145 0.0527417
R6178 VDD.n2148 VDD.n2147 0.0527417
R6179 VDD.n2150 VDD.n2149 0.0527417
R6180 VDD.n2152 VDD.n2151 0.0527417
R6181 VDD.n2154 VDD.n2153 0.0527417
R6182 VDD.n1939 VDD.n1938 0.0527417
R6183 VDD.n1941 VDD.n1940 0.0527417
R6184 VDD.n1943 VDD.n1942 0.0527417
R6185 VDD.n1945 VDD.n1944 0.0527417
R6186 VDD.n1947 VDD.n1946 0.0527417
R6187 VDD.n1949 VDD.n1948 0.0527417
R6188 VDD.n1951 VDD.n1950 0.0527417
R6189 VDD.n1953 VDD.n1952 0.0527417
R6190 VDD.n1955 VDD.n1954 0.0527417
R6191 VDD.n1957 VDD.n1956 0.0527417
R6192 VDD.n1959 VDD.n1958 0.0527417
R6193 VDD.n1961 VDD.n1960 0.0527417
R6194 VDD.n1963 VDD.n1962 0.0527417
R6195 VDD.n1965 VDD.n1964 0.0527417
R6196 VDD.n1967 VDD.n1966 0.0527417
R6197 VDD.n1969 VDD.n1968 0.0527417
R6198 VDD.n1971 VDD.n1970 0.0527417
R6199 VDD.n1973 VDD.n1972 0.0527417
R6200 VDD.n1975 VDD.n1974 0.0527417
R6201 VDD.n3057 VDD.n3056 0.0525833
R6202 VDD.n3061 VDD.n3060 0.0525833
R6203 VDD.n3065 VDD.n3064 0.0525833
R6204 VDD.n3088 VDD.n3087 0.0525833
R6205 VDD.n3092 VDD.n3091 0.0525833
R6206 VDD.n3096 VDD.n3095 0.0525833
R6207 VDD.n3119 VDD.n3118 0.0525833
R6208 VDD.n3123 VDD.n3122 0.0525833
R6209 VDD.n3127 VDD.n3126 0.0525833
R6210 VDD.n3150 VDD.n3149 0.0525833
R6211 VDD.n3154 VDD.n3153 0.0525833
R6212 VDD.n3158 VDD.n3157 0.0525833
R6213 VDD.n3181 VDD.n3180 0.0525833
R6214 VDD.n3185 VDD.n3184 0.0525833
R6215 VDD.n3189 VDD.n3188 0.0525833
R6216 VDD.n3212 VDD.n3211 0.0525833
R6217 VDD.n3216 VDD.n3215 0.0525833
R6218 VDD.n3220 VDD.n3219 0.0525833
R6219 VDD.n3243 VDD.n3242 0.0525833
R6220 VDD.n3247 VDD.n3246 0.0525833
R6221 VDD.n3251 VDD.n3250 0.0525833
R6222 VDD.n3274 VDD.n3273 0.0525833
R6223 VDD.n3278 VDD.n3277 0.0525833
R6224 VDD.n3282 VDD.n3281 0.0525833
R6225 VDD.n3305 VDD.n3304 0.0525833
R6226 VDD.n3309 VDD.n3308 0.0525833
R6227 VDD.n3313 VDD.n3312 0.0525833
R6228 VDD.n3336 VDD.n3335 0.0525833
R6229 VDD.n3340 VDD.n3339 0.0525833
R6230 VDD.n3344 VDD.n3343 0.0525833
R6231 VDD.n3367 VDD.n3366 0.0525833
R6232 VDD.n3371 VDD.n3370 0.0525833
R6233 VDD.n3375 VDD.n3374 0.0525833
R6234 VDD.n3024 VDD.n3023 0.0525833
R6235 VDD.n3408 VDD.n3407 0.0525833
R6236 VDD.n3428 VDD.n3427 0.0525833
R6237 VDD.n3448 VDD.n3447 0.0525833
R6238 VDD.n3469 VDD.n3468 0.0525833
R6239 VDD.n3536 VDD.n3534 0.0525833
R6240 VDD.n3579 VDD.n3578 0.0525833
R6241 VDD.n3599 VDD.n3598 0.0525833
R6242 VDD.n3619 VDD.n3618 0.0525833
R6243 VDD.n3639 VDD.n3638 0.0525833
R6244 VDD.n3712 VDD.n3709 0.0525833
R6245 VDD.n3750 VDD.n3749 0.0525833
R6246 VDD.n3770 VDD.n3769 0.0525833
R6247 VDD.n3789 VDD.n3788 0.0525833
R6248 VDD.n3810 VDD.n3809 0.0525833
R6249 VDD.n3888 VDD.n3886 0.0525833
R6250 VDD.n3918 VDD.n3917 0.0525833
R6251 VDD.n3938 VDD.n3937 0.0525833
R6252 VDD.n3958 VDD.n3957 0.0525833
R6253 VDD.n3979 VDD.n3978 0.0525833
R6254 VDD.n4085 VDD.n4084 0.0525833
R6255 VDD.n4103 VDD.n4102 0.0525833
R6256 VDD.n4121 VDD.n4120 0.0525833
R6257 VDD.n4140 VDD.n4139 0.0525833
R6258 VDD.n4232 VDD.n4231 0.0525833
R6259 VDD.n4252 VDD.n4251 0.0525833
R6260 VDD.n4270 VDD.n4269 0.0525833
R6261 VDD.n4289 VDD.n4288 0.0525833
R6262 VDD.n4388 VDD.n4387 0.0525833
R6263 VDD.n4406 VDD.n4405 0.0525833
R6264 VDD.n4424 VDD.n4423 0.0525833
R6265 VDD.n4443 VDD.n4442 0.0525833
R6266 VDD.n4525 VDD.n4510 0.0525833
R6267 VDD.n4551 VDD.n4550 0.0525833
R6268 VDD.n4560 VDD.n4559 0.0525833
R6269 VDD.n4584 VDD.n4583 0.0525833
R6270 VDD.n4605 VDD.n4604 0.0525833
R6271 VDD.n4677 VDD.n4675 0.0525833
R6272 VDD.n4716 VDD.n4715 0.0525833
R6273 VDD.n4735 VDD.n4734 0.0525833
R6274 VDD.n4755 VDD.n4754 0.0525833
R6275 VDD.n4772 VDD.n4771 0.0525833
R6276 VDD.n4846 VDD.n4842 0.0525833
R6277 VDD.n4881 VDD.n4880 0.0525833
R6278 VDD.n4905 VDD.n4904 0.0525833
R6279 VDD.n4914 VDD.n4913 0.0525833
R6280 VDD.n5011 VDD.n5009 0.0525833
R6281 VDD.n5050 VDD.n5049 0.0525833
R6282 VDD.n5070 VDD.n5069 0.0525833
R6283 VDD.n5088 VDD.n5087 0.0525833
R6284 VDD.n4353 VDD.n4351 0.0505
R6285 VDD.n4939 VDD.n4938 0.0505
R6286 VDD.n3047 VDD.n3046 0.0486358
R6287 VDD.n3071 VDD.n3070 0.0484167
R6288 VDD.n3075 VDD.n3074 0.0484167
R6289 VDD.n3079 VDD.n3078 0.0484167
R6290 VDD.n3102 VDD.n3101 0.0484167
R6291 VDD.n3106 VDD.n3105 0.0484167
R6292 VDD.n3110 VDD.n3109 0.0484167
R6293 VDD.n3133 VDD.n3132 0.0484167
R6294 VDD.n3137 VDD.n3136 0.0484167
R6295 VDD.n3141 VDD.n3140 0.0484167
R6296 VDD.n3164 VDD.n3163 0.0484167
R6297 VDD.n3168 VDD.n3167 0.0484167
R6298 VDD.n3172 VDD.n3171 0.0484167
R6299 VDD.n3195 VDD.n3194 0.0484167
R6300 VDD.n3199 VDD.n3198 0.0484167
R6301 VDD.n3203 VDD.n3202 0.0484167
R6302 VDD.n3226 VDD.n3225 0.0484167
R6303 VDD.n3230 VDD.n3229 0.0484167
R6304 VDD.n3234 VDD.n3233 0.0484167
R6305 VDD.n3257 VDD.n3256 0.0484167
R6306 VDD.n3261 VDD.n3260 0.0484167
R6307 VDD.n3265 VDD.n3264 0.0484167
R6308 VDD.n3288 VDD.n3287 0.0484167
R6309 VDD.n3292 VDD.n3291 0.0484167
R6310 VDD.n3296 VDD.n3295 0.0484167
R6311 VDD.n3319 VDD.n3318 0.0484167
R6312 VDD.n3323 VDD.n3322 0.0484167
R6313 VDD.n3327 VDD.n3326 0.0484167
R6314 VDD.n3350 VDD.n3349 0.0484167
R6315 VDD.n3354 VDD.n3353 0.0484167
R6316 VDD.n3358 VDD.n3357 0.0484167
R6317 VDD.n3381 VDD.n3380 0.0484167
R6318 VDD.n3385 VDD.n3384 0.0484167
R6319 VDD.n3389 VDD.n3388 0.0484167
R6320 VDD.n4215 VDD.n4203 0.0484167
R6321 VDD.n5107 VDD.n5106 0.0484167
R6322 VDD.n3047 VDD.n3001 0.048129
R6323 VDD.n4050 VDD.n4048 0.0463333
R6324 VDD.n3058 VDD.n3057 0.04425
R6325 VDD.n3060 VDD.n3059 0.04425
R6326 VDD.n3076 VDD.n3075 0.04425
R6327 VDD.n3078 VDD.n3077 0.04425
R6328 VDD.n3089 VDD.n3088 0.04425
R6329 VDD.n3091 VDD.n3090 0.04425
R6330 VDD.n3107 VDD.n3106 0.04425
R6331 VDD.n3109 VDD.n3108 0.04425
R6332 VDD.n3120 VDD.n3119 0.04425
R6333 VDD.n3122 VDD.n3121 0.04425
R6334 VDD.n3138 VDD.n3137 0.04425
R6335 VDD.n3140 VDD.n3139 0.04425
R6336 VDD.n3151 VDD.n3150 0.04425
R6337 VDD.n3153 VDD.n3152 0.04425
R6338 VDD.n3169 VDD.n3168 0.04425
R6339 VDD.n3171 VDD.n3170 0.04425
R6340 VDD.n3182 VDD.n3181 0.04425
R6341 VDD.n3184 VDD.n3183 0.04425
R6342 VDD.n3200 VDD.n3199 0.04425
R6343 VDD.n3202 VDD.n3201 0.04425
R6344 VDD.n3213 VDD.n3212 0.04425
R6345 VDD.n3215 VDD.n3214 0.04425
R6346 VDD.n3231 VDD.n3230 0.04425
R6347 VDD.n3233 VDD.n3232 0.04425
R6348 VDD.n3244 VDD.n3243 0.04425
R6349 VDD.n3246 VDD.n3245 0.04425
R6350 VDD.n3262 VDD.n3261 0.04425
R6351 VDD.n3264 VDD.n3263 0.04425
R6352 VDD.n3275 VDD.n3274 0.04425
R6353 VDD.n3277 VDD.n3276 0.04425
R6354 VDD.n3293 VDD.n3292 0.04425
R6355 VDD.n3295 VDD.n3294 0.04425
R6356 VDD.n3306 VDD.n3305 0.04425
R6357 VDD.n3308 VDD.n3307 0.04425
R6358 VDD.n3324 VDD.n3323 0.04425
R6359 VDD.n3326 VDD.n3325 0.04425
R6360 VDD.n3337 VDD.n3336 0.04425
R6361 VDD.n3339 VDD.n3338 0.04425
R6362 VDD.n3355 VDD.n3354 0.04425
R6363 VDD.n3357 VDD.n3356 0.04425
R6364 VDD.n3368 VDD.n3367 0.04425
R6365 VDD.n3370 VDD.n3369 0.04425
R6366 VDD.n3386 VDD.n3385 0.04425
R6367 VDD.n3388 VDD.n3387 0.04425
R6368 VDD.n3519 VDD.n3518 0.04425
R6369 VDD.n3525 VDD.n3520 0.04425
R6370 VDD.n3685 VDD.n3684 0.04425
R6371 VDD.n3856 VDD.n3855 0.04425
R6372 VDD.n3877 VDD.n3857 0.04425
R6373 VDD.n4025 VDD.n4024 0.04425
R6374 VDD.n4030 VDD.n4026 0.04425
R6375 VDD.n4181 VDD.n4180 0.04425
R6376 VDD.n4195 VDD.n4182 0.04425
R6377 VDD.n4329 VDD.n4328 0.04425
R6378 VDD.n4334 VDD.n4330 0.04425
R6379 VDD.n4486 VDD.n4485 0.04425
R6380 VDD.n4502 VDD.n4487 0.04425
R6381 VDD.n4557 VDD.n4551 0.04425
R6382 VDD.n4559 VDD.n4558 0.04425
R6383 VDD.n4651 VDD.n4650 0.04425
R6384 VDD.n4656 VDD.n4652 0.04425
R6385 VDD.n4734 VDD.n4733 0.04425
R6386 VDD.n4818 VDD.n4817 0.04425
R6387 VDD.n4836 VDD.n4819 0.04425
R6388 VDD.n4985 VDD.n4984 0.04425
R6389 VDD.n4990 VDD.n4986 0.04425
R6390 VDD.n5147 VDD.n5146 0.04425
R6391 VDD.n5152 VDD.n5148 0.04425
R6392 VDD.n3072 VDD.n3071 0.0421667
R6393 VDD.n3074 VDD.n3073 0.0421667
R6394 VDD.n3103 VDD.n3102 0.0421667
R6395 VDD.n3105 VDD.n3104 0.0421667
R6396 VDD.n3134 VDD.n3133 0.0421667
R6397 VDD.n3136 VDD.n3135 0.0421667
R6398 VDD.n3165 VDD.n3164 0.0421667
R6399 VDD.n3167 VDD.n3166 0.0421667
R6400 VDD.n3196 VDD.n3195 0.0421667
R6401 VDD.n3198 VDD.n3197 0.0421667
R6402 VDD.n3227 VDD.n3226 0.0421667
R6403 VDD.n3229 VDD.n3228 0.0421667
R6404 VDD.n3258 VDD.n3257 0.0421667
R6405 VDD.n3260 VDD.n3259 0.0421667
R6406 VDD.n3289 VDD.n3288 0.0421667
R6407 VDD.n3291 VDD.n3290 0.0421667
R6408 VDD.n3320 VDD.n3319 0.0421667
R6409 VDD.n3322 VDD.n3321 0.0421667
R6410 VDD.n3351 VDD.n3350 0.0421667
R6411 VDD.n3353 VDD.n3352 0.0421667
R6412 VDD.n3382 VDD.n3381 0.0421667
R6413 VDD.n3384 VDD.n3383 0.0421667
R6414 VDD.n3492 VDD.n3491 0.0421667
R6415 VDD.n3662 VDD.n3661 0.0421667
R6416 VDD.n3687 VDD.n3686 0.0421667
R6417 VDD.n3833 VDD.n3832 0.0421667
R6418 VDD.n4002 VDD.n4001 0.0421667
R6419 VDD.n4161 VDD.n4160 0.0421667
R6420 VDD.n4175 VDD.n4162 0.0421667
R6421 VDD.n4308 VDD.n4307 0.0421667
R6422 VDD.n4312 VDD.n4309 0.0421667
R6423 VDD.n4389 VDD.n4388 0.0421667
R6424 VDD.n4463 VDD.n4462 0.0421667
R6425 VDD.n4478 VDD.n4464 0.0421667
R6426 VDD.n4628 VDD.n4627 0.0421667
R6427 VDD.n4632 VDD.n4629 0.0421667
R6428 VDD.n4795 VDD.n4794 0.0421667
R6429 VDD.n4810 VDD.n4796 0.0421667
R6430 VDD.n4904 VDD.n4903 0.0421667
R6431 VDD.n4962 VDD.n4961 0.0421667
R6432 VDD.n4966 VDD.n4963 0.0421667
R6433 VDD.n5128 VDD.n5127 0.0421667
R6434 VDD.n5141 VDD.n5129 0.0421667
R6435 VDD.n1255 VDD.n1254 0.0415256
R6436 VDD.n158 VDD.n157 0.0410878
R6437 VDD.n4004 VDD.n4003 0.0400833
R6438 VDD.n4233 VDD.n4232 0.0400833
R6439 VDD.n5069 VDD.n5068 0.0400833
R6440 VDD.n6420 VDD.n6419 0.038709
R6441 VDD.n6314 VDD.n6313 0.038709
R6442 VDD.n3062 VDD.n3061 0.038
R6443 VDD.n3064 VDD.n3063 0.038
R6444 VDD.n3093 VDD.n3092 0.038
R6445 VDD.n3095 VDD.n3094 0.038
R6446 VDD.n3124 VDD.n3123 0.038
R6447 VDD.n3126 VDD.n3125 0.038
R6448 VDD.n3155 VDD.n3154 0.038
R6449 VDD.n3157 VDD.n3156 0.038
R6450 VDD.n3186 VDD.n3185 0.038
R6451 VDD.n3188 VDD.n3187 0.038
R6452 VDD.n3217 VDD.n3216 0.038
R6453 VDD.n3219 VDD.n3218 0.038
R6454 VDD.n3248 VDD.n3247 0.038
R6455 VDD.n3250 VDD.n3249 0.038
R6456 VDD.n3279 VDD.n3278 0.038
R6457 VDD.n3281 VDD.n3280 0.038
R6458 VDD.n3310 VDD.n3309 0.038
R6459 VDD.n3312 VDD.n3311 0.038
R6460 VDD.n3341 VDD.n3340 0.038
R6461 VDD.n3343 VDD.n3342 0.038
R6462 VDD.n3372 VDD.n3371 0.038
R6463 VDD.n3374 VDD.n3373 0.038
R6464 VDD.n3771 VDD.n3770 0.038
R6465 VDD.n3835 VDD.n3834 0.038
R6466 VDD.n3939 VDD.n3938 0.038
R6467 VDD.n4086 VDD.n4085 0.038
R6468 VDD.n4104 VDD.n4103 0.038
R6469 VDD.n4253 VDD.n4252 0.038
R6470 VDD.n4407 VDD.n4406 0.038
R6471 VDD.n4561 VDD.n4560 0.038
R6472 VDD.n4736 VDD.n4735 0.038
R6473 VDD.n4906 VDD.n4905 0.038
R6474 VDD.n4913 VDD.n4912 0.038
R6475 VDD.n99 VDD.n98 0.0364195
R6476 VDD.n3049 VDD.n3048 0.0359167
R6477 VDD.n3056 VDD.n3055 0.0359167
R6478 VDD.n3080 VDD.n3079 0.0359167
R6479 VDD.n3087 VDD.n3086 0.0359167
R6480 VDD.n3111 VDD.n3110 0.0359167
R6481 VDD.n3118 VDD.n3117 0.0359167
R6482 VDD.n3142 VDD.n3141 0.0359167
R6483 VDD.n3149 VDD.n3148 0.0359167
R6484 VDD.n3173 VDD.n3172 0.0359167
R6485 VDD.n3180 VDD.n3179 0.0359167
R6486 VDD.n3204 VDD.n3203 0.0359167
R6487 VDD.n3211 VDD.n3210 0.0359167
R6488 VDD.n3235 VDD.n3234 0.0359167
R6489 VDD.n3242 VDD.n3241 0.0359167
R6490 VDD.n3266 VDD.n3265 0.0359167
R6491 VDD.n3273 VDD.n3272 0.0359167
R6492 VDD.n3297 VDD.n3296 0.0359167
R6493 VDD.n3304 VDD.n3303 0.0359167
R6494 VDD.n3328 VDD.n3327 0.0359167
R6495 VDD.n3335 VDD.n3334 0.0359167
R6496 VDD.n3359 VDD.n3358 0.0359167
R6497 VDD.n3366 VDD.n3365 0.0359167
R6498 VDD.n5356 VDD.n3389 0.0359167
R6499 VDD.n3533 VDD.n3532 0.0359167
R6500 VDD.n3600 VDD.n3599 0.0359167
R6501 VDD.n3664 VDD.n3663 0.0359167
R6502 VDD.n3708 VDD.n3707 0.0359167
R6503 VDD.n3885 VDD.n3884 0.0359167
R6504 VDD.n3919 VDD.n3918 0.0359167
R6505 VDD.n4047 VDD.n4046 0.0359167
R6506 VDD.n4202 VDD.n4201 0.0359167
R6507 VDD.n4231 VDD.n4230 0.0359167
R6508 VDD.n4350 VDD.n4349 0.0359167
R6509 VDD.n4387 VDD.n4386 0.0359167
R6510 VDD.n4509 VDD.n4508 0.0359167
R6511 VDD.n4528 VDD.n4525 0.0359167
R6512 VDD.n4550 VDD.n4549 0.0359167
R6513 VDD.n4674 VDD.n4673 0.0359167
R6514 VDD.n4715 VDD.n4714 0.0359167
R6515 VDD.n4771 VDD.n4769 0.0359167
R6516 VDD.n4841 VDD.n4840 0.0359167
R6517 VDD.n4880 VDD.n4879 0.0359167
R6518 VDD.n5049 VDD.n5048 0.0359167
R6519 VDD.n5087 VDD.n5086 0.0359167
R6520 VDD.n3070 VDD.n3069 0.0338333
R6521 VDD.n3101 VDD.n3100 0.0338333
R6522 VDD.n3132 VDD.n3131 0.0338333
R6523 VDD.n3163 VDD.n3162 0.0338333
R6524 VDD.n3194 VDD.n3193 0.0338333
R6525 VDD.n3225 VDD.n3224 0.0338333
R6526 VDD.n3256 VDD.n3255 0.0338333
R6527 VDD.n3287 VDD.n3286 0.0338333
R6528 VDD.n3318 VDD.n3317 0.0338333
R6529 VDD.n3349 VDD.n3348 0.0338333
R6530 VDD.n3380 VDD.n3379 0.0338333
R6531 VDD.n3429 VDD.n3428 0.0338333
R6532 VDD.n3494 VDD.n3493 0.0338333
R6533 VDD.n3751 VDD.n3750 0.0338333
R6534 VDD.n4303 VDD.n4294 0.0338333
R6535 VDD.n4356 VDD.n4355 0.0338333
R6536 VDD.n4384 VDD.n4372 0.0338333
R6537 VDD.n4456 VDD.n4444 0.0338333
R6538 VDD.n4457 VDD.n4456 0.0338333
R6539 VDD.n4600 VDD.n4589 0.0338333
R6540 VDD.n4609 VDD.n4606 0.0338333
R6541 VDD.n4693 VDD.n4679 0.0338333
R6542 VDD.n4732 VDD.n4718 0.0338333
R6543 VDD.n4753 VDD.n4751 0.0338333
R6544 VDD.n4787 VDD.n4773 0.0338333
R6545 VDD.n4921 VDD.n4919 0.0338333
R6546 VDD.n4943 VDD.n4940 0.0338333
R6547 VDD.n5008 VDD.n5007 0.0338333
R6548 VDD.n5120 VDD.n5108 0.0338333
R6549 VDD.n3580 VDD.n3579 0.03175
R6550 VDD.n4155 VDD.n4154 0.03175
R6551 VDD.n4218 VDD.n4217 0.03175
R6552 VDD.n4291 VDD.n4290 0.03175
R6553 VDD.n4404 VDD.n4402 0.03175
R6554 VDD.n4440 VDD.n4438 0.03175
R6555 VDD.n4547 VDD.n4531 0.03175
R6556 VDD.n4582 VDD.n4565 0.03175
R6557 VDD.n4611 VDD.n4610 0.03175
R6558 VDD.n4840 VDD.n4838 0.03175
R6559 VDD.n4858 VDD.n4847 0.03175
R6560 VDD.n4901 VDD.n4882 0.03175
R6561 VDD.n5006 VDD.n4992 0.03175
R6562 VDD.n5104 VDD.n5102 0.03175
R6563 VDD.n5269 VDD.n5266 0.03175
R6564 VDD.n5355 VDD.n5270 0.03175
R6565 VDD.n111 VDD.n110 0.0302619
R6566 VDD.n3066 VDD.n3065 0.0296667
R6567 VDD.n3097 VDD.n3096 0.0296667
R6568 VDD.n3128 VDD.n3127 0.0296667
R6569 VDD.n3159 VDD.n3158 0.0296667
R6570 VDD.n3190 VDD.n3189 0.0296667
R6571 VDD.n3221 VDD.n3220 0.0296667
R6572 VDD.n3252 VDD.n3251 0.0296667
R6573 VDD.n3283 VDD.n3282 0.0296667
R6574 VDD.n3314 VDD.n3313 0.0296667
R6575 VDD.n3345 VDD.n3344 0.0296667
R6576 VDD.n3376 VDD.n3375 0.0296667
R6577 VDD.n3407 VDD.n3406 0.0296667
R6578 VDD.n3409 VDD.n3408 0.0296667
R6579 VDD.n3449 VDD.n3448 0.0296667
R6580 VDD.n3620 VDD.n3619 0.0296667
R6581 VDD.n3790 VDD.n3789 0.0296667
R6582 VDD.n3959 VDD.n3958 0.0296667
R6583 VDD.n3985 VDD.n3984 0.0296667
R6584 VDD.n4053 VDD.n4052 0.0296667
R6585 VDD.n4122 VDD.n4121 0.0296667
R6586 VDD.n4142 VDD.n4141 0.0296667
R6587 VDD.n4250 VDD.n4237 0.0296667
R6588 VDD.n4271 VDD.n4270 0.0296667
R6589 VDD.n4284 VDD.n4283 0.0296667
R6590 VDD.n4422 VDD.n4421 0.0296667
R6591 VDD.n4425 VDD.n4424 0.0296667
R6592 VDD.n4585 VDD.n4584 0.0296667
R6593 VDD.n4659 VDD.n4658 0.0296667
R6594 VDD.n4712 VDD.n4697 0.0296667
R6595 VDD.n4756 VDD.n4755 0.0296667
R6596 VDD.n4789 VDD.n4788 0.0296667
R6597 VDD.n4915 VDD.n4914 0.0296667
R6598 VDD.n5027 VDD.n5012 0.0296667
R6599 VDD.n5066 VDD.n5051 0.0296667
R6600 VDD.n5089 VDD.n5088 0.0296667
R6601 VDD.n901 VDD.n115 0.0294855
R6602 VDD.n133 VDD.n127 0.0294855
R6603 VDD.n891 VDD.n159 0.0294855
R6604 VDD.n98 VDD.n97 0.0292356
R6605 VDD.n100 VDD.n99 0.0277989
R6606 VDD.n3052 VDD.n3051 0.0275833
R6607 VDD.n3053 VDD.n3052 0.0275833
R6608 VDD.n3083 VDD.n3082 0.0275833
R6609 VDD.n3084 VDD.n3083 0.0275833
R6610 VDD.n3114 VDD.n3113 0.0275833
R6611 VDD.n3115 VDD.n3114 0.0275833
R6612 VDD.n3145 VDD.n3144 0.0275833
R6613 VDD.n3146 VDD.n3145 0.0275833
R6614 VDD.n3176 VDD.n3175 0.0275833
R6615 VDD.n3177 VDD.n3176 0.0275833
R6616 VDD.n3207 VDD.n3206 0.0275833
R6617 VDD.n3208 VDD.n3207 0.0275833
R6618 VDD.n3238 VDD.n3237 0.0275833
R6619 VDD.n3239 VDD.n3238 0.0275833
R6620 VDD.n3269 VDD.n3268 0.0275833
R6621 VDD.n3270 VDD.n3269 0.0275833
R6622 VDD.n3300 VDD.n3299 0.0275833
R6623 VDD.n3301 VDD.n3300 0.0275833
R6624 VDD.n3331 VDD.n3330 0.0275833
R6625 VDD.n3332 VDD.n3331 0.0275833
R6626 VDD.n3362 VDD.n3361 0.0275833
R6627 VDD.n3363 VDD.n3362 0.0275833
R6628 VDD.n3004 VDD.n3003 0.0275833
R6629 VDD.n3559 VDD.n3558 0.0275833
R6630 VDD.n3578 VDD.n3577 0.0275833
R6631 VDD.n3730 VDD.n3729 0.0275833
R6632 VDD.n3827 VDD.n3826 0.0275833
R6633 VDD.n3889 VDD.n3888 0.0275833
R6634 VDD.n3895 VDD.n3894 0.0275833
R6635 VDD.n3896 VDD.n3895 0.0275833
R6636 VDD.n3981 VDD.n3980 0.0275833
R6637 VDD.n4066 VDD.n4065 0.0275833
R6638 VDD.n4067 VDD.n4066 0.0275833
R6639 VDD.n4101 VDD.n4100 0.0275833
R6640 VDD.n4137 VDD.n4136 0.0275833
R6641 VDD.n4222 VDD.n4221 0.0275833
R6642 VDD.n4223 VDD.n4222 0.0275833
R6643 VDD.n4268 VDD.n4267 0.0275833
R6644 VDD.n4369 VDD.n4368 0.0275833
R6645 VDD.n4370 VDD.n4369 0.0275833
R6646 VDD.n4505 VDD.n4504 0.0275833
R6647 VDD.n4529 VDD.n4528 0.0275833
R6648 VDD.n4530 VDD.n4529 0.0275833
R6649 VDD.n4696 VDD.n4695 0.0275833
R6650 VDD.n4861 VDD.n4860 0.0275833
R6651 VDD.n4877 VDD.n4862 0.0275833
R6652 VDD.n4945 VDD.n4944 0.0275833
R6653 VDD.n5030 VDD.n5029 0.0275833
R6654 VDD.n891 VDD.n879 0.0258623
R6655 VDD.n3067 VDD.n3066 0.0255
R6656 VDD.n3098 VDD.n3097 0.0255
R6657 VDD.n3129 VDD.n3128 0.0255
R6658 VDD.n3160 VDD.n3159 0.0255
R6659 VDD.n3191 VDD.n3190 0.0255
R6660 VDD.n3222 VDD.n3221 0.0255
R6661 VDD.n3253 VDD.n3252 0.0255
R6662 VDD.n3284 VDD.n3283 0.0255
R6663 VDD.n3315 VDD.n3314 0.0255
R6664 VDD.n3346 VDD.n3345 0.0255
R6665 VDD.n3377 VDD.n3376 0.0255
R6666 VDD.n3427 VDD.n3426 0.0255
R6667 VDD.n3513 VDD.n3512 0.0255
R6668 VDD.n3645 VDD.n3644 0.0255
R6669 VDD.n3668 VDD.n3667 0.0255
R6670 VDD.n3713 VDD.n3712 0.0255
R6671 VDD.n3728 VDD.n3727 0.0255
R6672 VDD.n3749 VDD.n3748 0.0255
R6673 VDD.n3812 VDD.n3811 0.0255
R6674 VDD.n3850 VDD.n3849 0.0255
R6675 VDD.n3936 VDD.n3935 0.0255
R6676 VDD.n3974 VDD.n3973 0.0255
R6677 VDD.n4008 VDD.n4007 0.0255
R6678 VDD.n4119 VDD.n4118 0.0255
R6679 VDD.n4176 VDD.n4175 0.0255
R6680 VDD.n4337 VDD.n4336 0.0255
R6681 VDD.n4695 VDD.n4694 0.0255
R6682 VDD.n4769 VDD.n4756 0.0255
R6683 VDD.n4918 VDD.n4915 0.0255
R6684 VDD.n5046 VDD.n5031 0.0255
R6685 VDD.n5101 VDD.n5089 0.0255
R6686 VDD.n5122 VDD.n5121 0.0255
R6687 VDD.n902 VDD.n901 0.0249565
R6688 VDD VDD.n6709 0.0247117
R6689 VDD.n112 VDD.n111 0.0243095
R6690 VDD.n95 VDD.n92 0.0234885
R6691 VDD.n3487 VDD.n3486 0.0234167
R6692 VDD.n3537 VDD.n3536 0.0234167
R6693 VDD.n3557 VDD.n3556 0.0234167
R6694 VDD.n3598 VDD.n3597 0.0234167
R6695 VDD.n3641 VDD.n3640 0.0234167
R6696 VDD.n3768 VDD.n3767 0.0234167
R6697 VDD.n3807 VDD.n3806 0.0234167
R6698 VDD.n3917 VDD.n3916 0.0234167
R6699 VDD.n3956 VDD.n3955 0.0234167
R6700 VDD.n4198 VDD.n4197 0.0234167
R6701 VDD.n4314 VDD.n4313 0.0234167
R6702 VDD.n4586 VDD.n4585 0.0234167
R6703 VDD.n4860 VDD.n4859 0.0234167
R6704 VDD.n5146 VDD.n5143 0.0234167
R6705 VDD.n114 VDD.n113 0.023119
R6706 VDD.n110 VDD.n109 0.023119
R6707 VDD.n6213 VDD.n6212 0.0219844
R6708 VDD.n6206 VDD.n6205 0.0219844
R6709 VDD.n6199 VDD.n6198 0.0219844
R6710 VDD.n6192 VDD.n6191 0.0219844
R6711 VDD.n6185 VDD.n6184 0.0219844
R6712 VDD.n6178 VDD.n6177 0.0219844
R6713 VDD.n6171 VDD.n6170 0.0219844
R6714 VDD.n6164 VDD.n6163 0.0219844
R6715 VDD.n6157 VDD.n6156 0.0219844
R6716 VDD.n6150 VDD.n6149 0.0219844
R6717 VDD.n6143 VDD.n6142 0.0219844
R6718 VDD.n6136 VDD.n6135 0.0219844
R6719 VDD.n6129 VDD.n6128 0.0219844
R6720 VDD.n6122 VDD.n6121 0.0219844
R6721 VDD.n6115 VDD.n6114 0.0219844
R6722 VDD.n6108 VDD.n6107 0.0219844
R6723 VDD.n6101 VDD.n6100 0.0219844
R6724 VDD.n6094 VDD.n6093 0.0219844
R6725 VDD.n6087 VDD.n6086 0.0219844
R6726 VDD.n6080 VDD.n6079 0.0219844
R6727 VDD.n6034 VDD.n6033 0.0219844
R6728 VDD.n6027 VDD.n6026 0.0219844
R6729 VDD.n6020 VDD.n6019 0.0219844
R6730 VDD.n6013 VDD.n6012 0.0219844
R6731 VDD.n6006 VDD.n6005 0.0219844
R6732 VDD.n5999 VDD.n5998 0.0219844
R6733 VDD.n5992 VDD.n5991 0.0219844
R6734 VDD.n5985 VDD.n5984 0.0219844
R6735 VDD.n5978 VDD.n5977 0.0219844
R6736 VDD.n5971 VDD.n5970 0.0219844
R6737 VDD.n5964 VDD.n5963 0.0219844
R6738 VDD.n5957 VDD.n5956 0.0219844
R6739 VDD.n5950 VDD.n5949 0.0219844
R6740 VDD.n5943 VDD.n5942 0.0219844
R6741 VDD.n5936 VDD.n5935 0.0219844
R6742 VDD.n5929 VDD.n5928 0.0219844
R6743 VDD.n5922 VDD.n5921 0.0219844
R6744 VDD.n5915 VDD.n5914 0.0219844
R6745 VDD.n5908 VDD.n5907 0.0219844
R6746 VDD.n5901 VDD.n5900 0.0219844
R6747 VDD.n5855 VDD.n5854 0.0219844
R6748 VDD.n5848 VDD.n5847 0.0219844
R6749 VDD.n5841 VDD.n5840 0.0219844
R6750 VDD.n5834 VDD.n5833 0.0219844
R6751 VDD.n5827 VDD.n5826 0.0219844
R6752 VDD.n5820 VDD.n5819 0.0219844
R6753 VDD.n5813 VDD.n5812 0.0219844
R6754 VDD.n5806 VDD.n5805 0.0219844
R6755 VDD.n5799 VDD.n5798 0.0219844
R6756 VDD.n5792 VDD.n5791 0.0219844
R6757 VDD.n5785 VDD.n5784 0.0219844
R6758 VDD.n5778 VDD.n5777 0.0219844
R6759 VDD.n5771 VDD.n5770 0.0219844
R6760 VDD.n5764 VDD.n5763 0.0219844
R6761 VDD.n5757 VDD.n5756 0.0219844
R6762 VDD.n5750 VDD.n5749 0.0219844
R6763 VDD.n5743 VDD.n5742 0.0219844
R6764 VDD.n5736 VDD.n5735 0.0219844
R6765 VDD.n5729 VDD.n5728 0.0219844
R6766 VDD.n5722 VDD.n5721 0.0219844
R6767 VDD.n5676 VDD.n5675 0.0219844
R6768 VDD.n5669 VDD.n5668 0.0219844
R6769 VDD.n5662 VDD.n5661 0.0219844
R6770 VDD.n5655 VDD.n5654 0.0219844
R6771 VDD.n5648 VDD.n5647 0.0219844
R6772 VDD.n5641 VDD.n5640 0.0219844
R6773 VDD.n5634 VDD.n5633 0.0219844
R6774 VDD.n5627 VDD.n5626 0.0219844
R6775 VDD.n5620 VDD.n5619 0.0219844
R6776 VDD.n5613 VDD.n5612 0.0219844
R6777 VDD.n5606 VDD.n5605 0.0219844
R6778 VDD.n5599 VDD.n5598 0.0219844
R6779 VDD.n5592 VDD.n5591 0.0219844
R6780 VDD.n5585 VDD.n5584 0.0219844
R6781 VDD.n5578 VDD.n5577 0.0219844
R6782 VDD.n5571 VDD.n5570 0.0219844
R6783 VDD.n5564 VDD.n5563 0.0219844
R6784 VDD.n5557 VDD.n5556 0.0219844
R6785 VDD.n5550 VDD.n5549 0.0219844
R6786 VDD.n5543 VDD.n5542 0.0219844
R6787 VDD.n5497 VDD.n5496 0.0219844
R6788 VDD.n5490 VDD.n5489 0.0219844
R6789 VDD.n5483 VDD.n5482 0.0219844
R6790 VDD.n5476 VDD.n5475 0.0219844
R6791 VDD.n5469 VDD.n5468 0.0219844
R6792 VDD.n5462 VDD.n5461 0.0219844
R6793 VDD.n5455 VDD.n5454 0.0219844
R6794 VDD.n5448 VDD.n5447 0.0219844
R6795 VDD.n5441 VDD.n5440 0.0219844
R6796 VDD.n5434 VDD.n5433 0.0219844
R6797 VDD.n5427 VDD.n5426 0.0219844
R6798 VDD.n5420 VDD.n5419 0.0219844
R6799 VDD.n5413 VDD.n5412 0.0219844
R6800 VDD.n5406 VDD.n5405 0.0219844
R6801 VDD.n5399 VDD.n5398 0.0219844
R6802 VDD.n5392 VDD.n5391 0.0219844
R6803 VDD.n5385 VDD.n5384 0.0219844
R6804 VDD.n5378 VDD.n5377 0.0219844
R6805 VDD.n5371 VDD.n5370 0.0219844
R6806 VDD.n5364 VDD.n5363 0.0219844
R6807 VDD.n2652 VDD.n2651 0.0219844
R6808 VDD.n2645 VDD.n2644 0.0219844
R6809 VDD.n2638 VDD.n2637 0.0219844
R6810 VDD.n2631 VDD.n2630 0.0219844
R6811 VDD.n2624 VDD.n2623 0.0219844
R6812 VDD.n2617 VDD.n2616 0.0219844
R6813 VDD.n2610 VDD.n2609 0.0219844
R6814 VDD.n2603 VDD.n2602 0.0219844
R6815 VDD.n2596 VDD.n2595 0.0219844
R6816 VDD.n2589 VDD.n2588 0.0219844
R6817 VDD.n2582 VDD.n2581 0.0219844
R6818 VDD.n2575 VDD.n2574 0.0219844
R6819 VDD.n2568 VDD.n2567 0.0219844
R6820 VDD.n2561 VDD.n2560 0.0219844
R6821 VDD.n2554 VDD.n2553 0.0219844
R6822 VDD.n2547 VDD.n2546 0.0219844
R6823 VDD.n2540 VDD.n2539 0.0219844
R6824 VDD.n2533 VDD.n2532 0.0219844
R6825 VDD.n2526 VDD.n2525 0.0219844
R6826 VDD.n2519 VDD.n2518 0.0219844
R6827 VDD.n2473 VDD.n2472 0.0219844
R6828 VDD.n2466 VDD.n2465 0.0219844
R6829 VDD.n2459 VDD.n2458 0.0219844
R6830 VDD.n2452 VDD.n2451 0.0219844
R6831 VDD.n2445 VDD.n2444 0.0219844
R6832 VDD.n2438 VDD.n2437 0.0219844
R6833 VDD.n2431 VDD.n2430 0.0219844
R6834 VDD.n2424 VDD.n2423 0.0219844
R6835 VDD.n2417 VDD.n2416 0.0219844
R6836 VDD.n2410 VDD.n2409 0.0219844
R6837 VDD.n2403 VDD.n2402 0.0219844
R6838 VDD.n2396 VDD.n2395 0.0219844
R6839 VDD.n2389 VDD.n2388 0.0219844
R6840 VDD.n2382 VDD.n2381 0.0219844
R6841 VDD.n2375 VDD.n2374 0.0219844
R6842 VDD.n2368 VDD.n2367 0.0219844
R6843 VDD.n2361 VDD.n2360 0.0219844
R6844 VDD.n2354 VDD.n2353 0.0219844
R6845 VDD.n2347 VDD.n2346 0.0219844
R6846 VDD.n2340 VDD.n2339 0.0219844
R6847 VDD.n2294 VDD.n2293 0.0219844
R6848 VDD.n2287 VDD.n2286 0.0219844
R6849 VDD.n2280 VDD.n2279 0.0219844
R6850 VDD.n2273 VDD.n2272 0.0219844
R6851 VDD.n2266 VDD.n2265 0.0219844
R6852 VDD.n2259 VDD.n2258 0.0219844
R6853 VDD.n2252 VDD.n2251 0.0219844
R6854 VDD.n2245 VDD.n2244 0.0219844
R6855 VDD.n2238 VDD.n2237 0.0219844
R6856 VDD.n2231 VDD.n2230 0.0219844
R6857 VDD.n2224 VDD.n2223 0.0219844
R6858 VDD.n2217 VDD.n2216 0.0219844
R6859 VDD.n2210 VDD.n2209 0.0219844
R6860 VDD.n2203 VDD.n2202 0.0219844
R6861 VDD.n2196 VDD.n2195 0.0219844
R6862 VDD.n2189 VDD.n2188 0.0219844
R6863 VDD.n2182 VDD.n2181 0.0219844
R6864 VDD.n2175 VDD.n2174 0.0219844
R6865 VDD.n2168 VDD.n2167 0.0219844
R6866 VDD.n2161 VDD.n2160 0.0219844
R6867 VDD.n2115 VDD.n2114 0.0219844
R6868 VDD.n2108 VDD.n2107 0.0219844
R6869 VDD.n2101 VDD.n2100 0.0219844
R6870 VDD.n2094 VDD.n2093 0.0219844
R6871 VDD.n2087 VDD.n2086 0.0219844
R6872 VDD.n2080 VDD.n2079 0.0219844
R6873 VDD.n2073 VDD.n2072 0.0219844
R6874 VDD.n2066 VDD.n2065 0.0219844
R6875 VDD.n2059 VDD.n2058 0.0219844
R6876 VDD.n2052 VDD.n2051 0.0219844
R6877 VDD.n2045 VDD.n2044 0.0219844
R6878 VDD.n2038 VDD.n2037 0.0219844
R6879 VDD.n2031 VDD.n2030 0.0219844
R6880 VDD.n2024 VDD.n2023 0.0219844
R6881 VDD.n2017 VDD.n2016 0.0219844
R6882 VDD.n2010 VDD.n2009 0.0219844
R6883 VDD.n2003 VDD.n2002 0.0219844
R6884 VDD.n1996 VDD.n1995 0.0219844
R6885 VDD.n1989 VDD.n1988 0.0219844
R6886 VDD.n1982 VDD.n1981 0.0219844
R6887 VDD.n1936 VDD.n1935 0.0219844
R6888 VDD.n1929 VDD.n1928 0.0219844
R6889 VDD.n1922 VDD.n1921 0.0219844
R6890 VDD.n1915 VDD.n1914 0.0219844
R6891 VDD.n1908 VDD.n1907 0.0219844
R6892 VDD.n1901 VDD.n1900 0.0219844
R6893 VDD.n1894 VDD.n1893 0.0219844
R6894 VDD.n1887 VDD.n1886 0.0219844
R6895 VDD.n1880 VDD.n1879 0.0219844
R6896 VDD.n1873 VDD.n1872 0.0219844
R6897 VDD.n1866 VDD.n1865 0.0219844
R6898 VDD.n1859 VDD.n1858 0.0219844
R6899 VDD.n1852 VDD.n1851 0.0219844
R6900 VDD.n1845 VDD.n1844 0.0219844
R6901 VDD.n1838 VDD.n1837 0.0219844
R6902 VDD.n1831 VDD.n1830 0.0219844
R6903 VDD.n1824 VDD.n1823 0.0219844
R6904 VDD.n1817 VDD.n1816 0.0219844
R6905 VDD.n1810 VDD.n1809 0.0219844
R6906 VDD.n1803 VDD.n1802 0.0219844
R6907 VDD.n3069 VDD.n3068 0.0213333
R6908 VDD.n3100 VDD.n3099 0.0213333
R6909 VDD.n3131 VDD.n3130 0.0213333
R6910 VDD.n3162 VDD.n3161 0.0213333
R6911 VDD.n3193 VDD.n3192 0.0213333
R6912 VDD.n3224 VDD.n3223 0.0213333
R6913 VDD.n3255 VDD.n3254 0.0213333
R6914 VDD.n3286 VDD.n3285 0.0213333
R6915 VDD.n3317 VDD.n3316 0.0213333
R6916 VDD.n3348 VDD.n3347 0.0213333
R6917 VDD.n3379 VDD.n3378 0.0213333
R6918 VDD.n3023 VDD.n3020 0.0213333
R6919 VDD.n3019 VDD.n3005 0.0213333
R6920 VDD.n3447 VDD.n3446 0.0213333
R6921 VDD.n3470 VDD.n3469 0.0213333
R6922 VDD.n3471 VDD.n3470 0.0213333
R6923 VDD.n3518 VDD.n3514 0.0213333
R6924 VDD.n3597 VDD.n3596 0.0213333
R6925 VDD.n3635 VDD.n3634 0.0213333
R6926 VDD.n3640 VDD.n3639 0.0213333
R6927 VDD.n3769 VDD.n3768 0.0213333
R6928 VDD.n3787 VDD.n3786 0.0213333
R6929 VDD.n3811 VDD.n3810 0.0213333
R6930 VDD.n3980 VDD.n3979 0.0213333
R6931 VDD.n4033 VDD.n4032 0.0213333
R6932 VDD.n4084 VDD.n4083 0.0213333
R6933 VDD.n4141 VDD.n4140 0.0213333
R6934 VDD.n4290 VDD.n4289 0.0213333
R6935 VDD.n4426 VDD.n4425 0.0213333
R6936 VDD.n4444 VDD.n4443 0.0213333
R6937 VDD.n4480 VDD.n4479 0.0213333
R6938 VDD.n4606 VDD.n4605 0.0213333
R6939 VDD.n4773 VDD.n4772 0.0213333
R6940 VDD.n4940 VDD.n4939 0.0213333
R6941 VDD.n4969 VDD.n4968 0.0213333
R6942 VDD.n5029 VDD.n5028 0.0213333
R6943 VDD.n5108 VDD.n5107 0.0213333
R6944 VDD.n148 VDD.n147 0.0208126
R6945 VDD.n140 VDD.n139 0.0203238
R6946 VDD.n142 VDD.n140 0.0203238
R6947 VDD.n153 VDD.n152 0.0203238
R6948 VDD.n152 VDD.n151 0.0203238
R6949 VDD.n151 VDD.n150 0.0203238
R6950 VDD.n150 VDD.n149 0.0203238
R6951 VDD.n149 VDD.n148 0.0203238
R6952 VDD.n3050 VDD.n3049 0.01925
R6953 VDD.n3055 VDD.n3054 0.01925
R6954 VDD.n3081 VDD.n3080 0.01925
R6955 VDD.n3086 VDD.n3085 0.01925
R6956 VDD.n3112 VDD.n3111 0.01925
R6957 VDD.n3117 VDD.n3116 0.01925
R6958 VDD.n3143 VDD.n3142 0.01925
R6959 VDD.n3148 VDD.n3147 0.01925
R6960 VDD.n3174 VDD.n3173 0.01925
R6961 VDD.n3179 VDD.n3178 0.01925
R6962 VDD.n3205 VDD.n3204 0.01925
R6963 VDD.n3210 VDD.n3209 0.01925
R6964 VDD.n3236 VDD.n3235 0.01925
R6965 VDD.n3241 VDD.n3240 0.01925
R6966 VDD.n3267 VDD.n3266 0.01925
R6967 VDD.n3272 VDD.n3271 0.01925
R6968 VDD.n3298 VDD.n3297 0.01925
R6969 VDD.n3303 VDD.n3302 0.01925
R6970 VDD.n3329 VDD.n3328 0.01925
R6971 VDD.n3334 VDD.n3333 0.01925
R6972 VDD.n3360 VDD.n3359 0.01925
R6973 VDD.n3365 VDD.n3364 0.01925
R6974 VDD.n5357 VDD.n5356 0.01925
R6975 VDD.n3041 VDD.n3040 0.01925
R6976 VDD.n3026 VDD.n3025 0.01925
R6977 VDD.n3025 VDD.n3024 0.01925
R6978 VDD.n3405 VDD.n3404 0.01925
R6979 VDD.n3426 VDD.n3425 0.01925
R6980 VDD.n3466 VDD.n3465 0.01925
R6981 VDD.n3534 VDD.n3533 0.01925
R6982 VDD.n3576 VDD.n3575 0.01925
R6983 VDD.n3617 VDD.n3616 0.01925
R6984 VDD.n3618 VDD.n3617 0.01925
R6985 VDD.n3684 VDD.n3669 0.01925
R6986 VDD.n3709 VDD.n3708 0.01925
R6987 VDD.n3747 VDD.n3746 0.01925
R6988 VDD.n3879 VDD.n3878 0.01925
R6989 VDD.n3886 VDD.n3885 0.01925
R6990 VDD.n3901 VDD.n3900 0.01925
R6991 VDD.n3937 VDD.n3936 0.01925
R6992 VDD.n4048 VDD.n4047 0.01925
R6993 VDD.n4081 VDD.n4080 0.01925
R6994 VDD.n4203 VDD.n4202 0.01925
R6995 VDD.n4230 VDD.n4229 0.01925
R6996 VDD.n4272 VDD.n4271 0.01925
R6997 VDD.n4351 VDD.n4350 0.01925
R6998 VDD.n4510 VDD.n4509 0.01925
R6999 VDD.n4634 VDD.n4633 0.01925
R7000 VDD.n4675 VDD.n4674 0.01925
R7001 VDD.n4813 VDD.n4812 0.01925
R7002 VDD.n4842 VDD.n4841 0.01925
R7003 VDD.n5009 VDD.n5008 0.01925
R7004 VDD.n5072 VDD.n5070 0.01925
R7005 VDD.n5073 VDD.n5072 0.01925
R7006 VDD.n5355 VDD.n5354 0.01925
R7007 VDD.n6212 VDD.n6209 0.0174092
R7008 VDD.n6205 VDD.n6202 0.0174092
R7009 VDD.n6198 VDD.n6195 0.0174092
R7010 VDD.n6191 VDD.n6188 0.0174092
R7011 VDD.n6184 VDD.n6181 0.0174092
R7012 VDD.n6177 VDD.n6174 0.0174092
R7013 VDD.n6170 VDD.n6167 0.0174092
R7014 VDD.n6163 VDD.n6160 0.0174092
R7015 VDD.n6156 VDD.n6153 0.0174092
R7016 VDD.n6149 VDD.n6146 0.0174092
R7017 VDD.n6142 VDD.n6139 0.0174092
R7018 VDD.n6135 VDD.n6132 0.0174092
R7019 VDD.n6128 VDD.n6125 0.0174092
R7020 VDD.n6121 VDD.n6118 0.0174092
R7021 VDD.n6114 VDD.n6111 0.0174092
R7022 VDD.n6107 VDD.n6104 0.0174092
R7023 VDD.n6100 VDD.n6097 0.0174092
R7024 VDD.n6093 VDD.n6090 0.0174092
R7025 VDD.n6086 VDD.n6083 0.0174092
R7026 VDD.n6079 VDD.n6076 0.0174092
R7027 VDD.n6033 VDD.n6030 0.0174092
R7028 VDD.n6026 VDD.n6023 0.0174092
R7029 VDD.n6019 VDD.n6016 0.0174092
R7030 VDD.n6012 VDD.n6009 0.0174092
R7031 VDD.n6005 VDD.n6002 0.0174092
R7032 VDD.n5998 VDD.n5995 0.0174092
R7033 VDD.n5991 VDD.n5988 0.0174092
R7034 VDD.n5984 VDD.n5981 0.0174092
R7035 VDD.n5977 VDD.n5974 0.0174092
R7036 VDD.n5970 VDD.n5967 0.0174092
R7037 VDD.n5963 VDD.n5960 0.0174092
R7038 VDD.n5956 VDD.n5953 0.0174092
R7039 VDD.n5949 VDD.n5946 0.0174092
R7040 VDD.n5942 VDD.n5939 0.0174092
R7041 VDD.n5935 VDD.n5932 0.0174092
R7042 VDD.n5928 VDD.n5925 0.0174092
R7043 VDD.n5921 VDD.n5918 0.0174092
R7044 VDD.n5914 VDD.n5911 0.0174092
R7045 VDD.n5907 VDD.n5904 0.0174092
R7046 VDD.n5900 VDD.n5897 0.0174092
R7047 VDD.n5854 VDD.n5851 0.0174092
R7048 VDD.n5847 VDD.n5844 0.0174092
R7049 VDD.n5840 VDD.n5837 0.0174092
R7050 VDD.n5833 VDD.n5830 0.0174092
R7051 VDD.n5826 VDD.n5823 0.0174092
R7052 VDD.n5819 VDD.n5816 0.0174092
R7053 VDD.n5812 VDD.n5809 0.0174092
R7054 VDD.n5805 VDD.n5802 0.0174092
R7055 VDD.n5798 VDD.n5795 0.0174092
R7056 VDD.n5791 VDD.n5788 0.0174092
R7057 VDD.n5784 VDD.n5781 0.0174092
R7058 VDD.n5777 VDD.n5774 0.0174092
R7059 VDD.n5770 VDD.n5767 0.0174092
R7060 VDD.n5763 VDD.n5760 0.0174092
R7061 VDD.n5756 VDD.n5753 0.0174092
R7062 VDD.n5749 VDD.n5746 0.0174092
R7063 VDD.n5742 VDD.n5739 0.0174092
R7064 VDD.n5735 VDD.n5732 0.0174092
R7065 VDD.n5728 VDD.n5725 0.0174092
R7066 VDD.n5721 VDD.n5718 0.0174092
R7067 VDD.n5675 VDD.n5672 0.0174092
R7068 VDD.n5668 VDD.n5665 0.0174092
R7069 VDD.n5661 VDD.n5658 0.0174092
R7070 VDD.n5654 VDD.n5651 0.0174092
R7071 VDD.n5647 VDD.n5644 0.0174092
R7072 VDD.n5640 VDD.n5637 0.0174092
R7073 VDD.n5633 VDD.n5630 0.0174092
R7074 VDD.n5626 VDD.n5623 0.0174092
R7075 VDD.n5619 VDD.n5616 0.0174092
R7076 VDD.n5612 VDD.n5609 0.0174092
R7077 VDD.n5605 VDD.n5602 0.0174092
R7078 VDD.n5598 VDD.n5595 0.0174092
R7079 VDD.n5591 VDD.n5588 0.0174092
R7080 VDD.n5584 VDD.n5581 0.0174092
R7081 VDD.n5577 VDD.n5574 0.0174092
R7082 VDD.n5570 VDD.n5567 0.0174092
R7083 VDD.n5563 VDD.n5560 0.0174092
R7084 VDD.n5556 VDD.n5553 0.0174092
R7085 VDD.n5549 VDD.n5546 0.0174092
R7086 VDD.n5542 VDD.n5539 0.0174092
R7087 VDD.n5496 VDD.n5493 0.0174092
R7088 VDD.n5489 VDD.n5486 0.0174092
R7089 VDD.n5482 VDD.n5479 0.0174092
R7090 VDD.n5475 VDD.n5472 0.0174092
R7091 VDD.n5468 VDD.n5465 0.0174092
R7092 VDD.n5461 VDD.n5458 0.0174092
R7093 VDD.n5454 VDD.n5451 0.0174092
R7094 VDD.n5447 VDD.n5444 0.0174092
R7095 VDD.n5440 VDD.n5437 0.0174092
R7096 VDD.n5433 VDD.n5430 0.0174092
R7097 VDD.n5426 VDD.n5423 0.0174092
R7098 VDD.n5419 VDD.n5416 0.0174092
R7099 VDD.n5412 VDD.n5409 0.0174092
R7100 VDD.n5405 VDD.n5402 0.0174092
R7101 VDD.n5398 VDD.n5395 0.0174092
R7102 VDD.n5391 VDD.n5388 0.0174092
R7103 VDD.n5384 VDD.n5381 0.0174092
R7104 VDD.n5377 VDD.n5374 0.0174092
R7105 VDD.n5370 VDD.n5367 0.0174092
R7106 VDD.n5363 VDD.n5360 0.0174092
R7107 VDD.n2651 VDD.n2650 0.0174092
R7108 VDD.n2644 VDD.n2643 0.0174092
R7109 VDD.n2637 VDD.n2636 0.0174092
R7110 VDD.n2630 VDD.n2629 0.0174092
R7111 VDD.n2623 VDD.n2622 0.0174092
R7112 VDD.n2616 VDD.n2615 0.0174092
R7113 VDD.n2609 VDD.n2608 0.0174092
R7114 VDD.n2602 VDD.n2601 0.0174092
R7115 VDD.n2595 VDD.n2594 0.0174092
R7116 VDD.n2588 VDD.n2587 0.0174092
R7117 VDD.n2581 VDD.n2580 0.0174092
R7118 VDD.n2574 VDD.n2573 0.0174092
R7119 VDD.n2567 VDD.n2566 0.0174092
R7120 VDD.n2560 VDD.n2559 0.0174092
R7121 VDD.n2553 VDD.n2552 0.0174092
R7122 VDD.n2546 VDD.n2545 0.0174092
R7123 VDD.n2539 VDD.n2538 0.0174092
R7124 VDD.n2532 VDD.n2531 0.0174092
R7125 VDD.n2525 VDD.n2524 0.0174092
R7126 VDD.n2518 VDD.n2517 0.0174092
R7127 VDD.n2472 VDD.n2471 0.0174092
R7128 VDD.n2465 VDD.n2464 0.0174092
R7129 VDD.n2458 VDD.n2457 0.0174092
R7130 VDD.n2451 VDD.n2450 0.0174092
R7131 VDD.n2444 VDD.n2443 0.0174092
R7132 VDD.n2437 VDD.n2436 0.0174092
R7133 VDD.n2430 VDD.n2429 0.0174092
R7134 VDD.n2423 VDD.n2422 0.0174092
R7135 VDD.n2416 VDD.n2415 0.0174092
R7136 VDD.n2409 VDD.n2408 0.0174092
R7137 VDD.n2402 VDD.n2401 0.0174092
R7138 VDD.n2395 VDD.n2394 0.0174092
R7139 VDD.n2388 VDD.n2387 0.0174092
R7140 VDD.n2381 VDD.n2380 0.0174092
R7141 VDD.n2374 VDD.n2373 0.0174092
R7142 VDD.n2367 VDD.n2366 0.0174092
R7143 VDD.n2360 VDD.n2359 0.0174092
R7144 VDD.n2353 VDD.n2352 0.0174092
R7145 VDD.n2346 VDD.n2345 0.0174092
R7146 VDD.n2339 VDD.n2338 0.0174092
R7147 VDD.n2293 VDD.n2292 0.0174092
R7148 VDD.n2286 VDD.n2285 0.0174092
R7149 VDD.n2279 VDD.n2278 0.0174092
R7150 VDD.n2272 VDD.n2271 0.0174092
R7151 VDD.n2265 VDD.n2264 0.0174092
R7152 VDD.n2258 VDD.n2257 0.0174092
R7153 VDD.n2251 VDD.n2250 0.0174092
R7154 VDD.n2244 VDD.n2243 0.0174092
R7155 VDD.n2237 VDD.n2236 0.0174092
R7156 VDD.n2230 VDD.n2229 0.0174092
R7157 VDD.n2223 VDD.n2222 0.0174092
R7158 VDD.n2216 VDD.n2215 0.0174092
R7159 VDD.n2209 VDD.n2208 0.0174092
R7160 VDD.n2202 VDD.n2201 0.0174092
R7161 VDD.n2195 VDD.n2194 0.0174092
R7162 VDD.n2188 VDD.n2187 0.0174092
R7163 VDD.n2181 VDD.n2180 0.0174092
R7164 VDD.n2174 VDD.n2173 0.0174092
R7165 VDD.n2167 VDD.n2166 0.0174092
R7166 VDD.n2160 VDD.n2159 0.0174092
R7167 VDD.n2114 VDD.n2111 0.0174092
R7168 VDD.n2107 VDD.n2104 0.0174092
R7169 VDD.n2100 VDD.n2097 0.0174092
R7170 VDD.n2093 VDD.n2090 0.0174092
R7171 VDD.n2086 VDD.n2083 0.0174092
R7172 VDD.n2079 VDD.n2076 0.0174092
R7173 VDD.n2072 VDD.n2069 0.0174092
R7174 VDD.n2065 VDD.n2062 0.0174092
R7175 VDD.n2058 VDD.n2055 0.0174092
R7176 VDD.n2051 VDD.n2048 0.0174092
R7177 VDD.n2044 VDD.n2041 0.0174092
R7178 VDD.n2037 VDD.n2034 0.0174092
R7179 VDD.n2030 VDD.n2027 0.0174092
R7180 VDD.n2023 VDD.n2020 0.0174092
R7181 VDD.n2016 VDD.n2013 0.0174092
R7182 VDD.n2009 VDD.n2006 0.0174092
R7183 VDD.n2002 VDD.n1999 0.0174092
R7184 VDD.n1995 VDD.n1992 0.0174092
R7185 VDD.n1988 VDD.n1985 0.0174092
R7186 VDD.n1981 VDD.n1978 0.0174092
R7187 VDD.n1935 VDD.n1932 0.0174092
R7188 VDD.n1928 VDD.n1925 0.0174092
R7189 VDD.n1921 VDD.n1918 0.0174092
R7190 VDD.n1914 VDD.n1911 0.0174092
R7191 VDD.n1907 VDD.n1904 0.0174092
R7192 VDD.n1900 VDD.n1897 0.0174092
R7193 VDD.n1893 VDD.n1890 0.0174092
R7194 VDD.n1886 VDD.n1883 0.0174092
R7195 VDD.n1879 VDD.n1876 0.0174092
R7196 VDD.n1872 VDD.n1869 0.0174092
R7197 VDD.n1865 VDD.n1862 0.0174092
R7198 VDD.n1858 VDD.n1855 0.0174092
R7199 VDD.n1851 VDD.n1848 0.0174092
R7200 VDD.n1844 VDD.n1841 0.0174092
R7201 VDD.n1837 VDD.n1834 0.0174092
R7202 VDD.n1830 VDD.n1827 0.0174092
R7203 VDD.n1823 VDD.n1820 0.0174092
R7204 VDD.n1816 VDD.n1813 0.0174092
R7205 VDD.n1809 VDD.n1806 0.0174092
R7206 VDD.n1802 VDD.n1799 0.0174092
R7207 VDD.n3046 VDD.n3042 0.0171667
R7208 VDD.n3040 VDD.n3026 0.0171667
R7209 VDD.n3446 VDD.n3445 0.0171667
R7210 VDD.n3465 VDD.n3450 0.0171667
R7211 VDD.n3468 VDD.n3466 0.0171667
R7212 VDD.n3526 VDD.n3525 0.0171667
R7213 VDD.n3532 VDD.n3527 0.0171667
R7214 VDD.n3692 VDD.n3691 0.0171667
R7215 VDD.n3693 VDD.n3692 0.0171667
R7216 VDD.n3788 VDD.n3787 0.0171667
R7217 VDD.n3855 VDD.n3851 0.0171667
R7218 VDD.n3878 VDD.n3877 0.0171667
R7219 VDD.n4102 VDD.n4101 0.0171667
R7220 VDD.n4123 VDD.n4122 0.0171667
R7221 VDD.n4386 VDD.n4385 0.0171667
R7222 VDD.n4635 VDD.n4634 0.0171667
R7223 VDD.n4812 VDD.n4811 0.0171667
R7224 VDD.n5266 VDD.n5152 0.0171667
R7225 VDD.n157 VDD.n156 0.0171052
R7226 VDD.n138 VDD.n137 0.0171052
R7227 VDD.n137 VDD.n136 0.0171052
R7228 VDD.n136 VDD.n135 0.0171052
R7229 VDD.n135 VDD.n134 0.0171052
R7230 VDD.n3063 VDD.n3062 0.0150833
R7231 VDD.n3094 VDD.n3093 0.0150833
R7232 VDD.n3125 VDD.n3124 0.0150833
R7233 VDD.n3156 VDD.n3155 0.0150833
R7234 VDD.n3187 VDD.n3186 0.0150833
R7235 VDD.n3218 VDD.n3217 0.0150833
R7236 VDD.n3249 VDD.n3248 0.0150833
R7237 VDD.n3280 VDD.n3279 0.0150833
R7238 VDD.n3311 VDD.n3310 0.0150833
R7239 VDD.n3342 VDD.n3341 0.0150833
R7240 VDD.n3373 VDD.n3372 0.0150833
R7241 VDD.n3020 VDD.n3019 0.0150833
R7242 VDD.n3424 VDD.n3409 0.0150833
R7243 VDD.n3445 VDD.n3430 0.0150833
R7244 VDD.n3491 VDD.n3488 0.0150833
R7245 VDD.n3527 VDD.n3526 0.0150833
R7246 VDD.n3616 VDD.n3601 0.0150833
R7247 VDD.n3634 VDD.n3621 0.0150833
R7248 VDD.n3638 VDD.n3635 0.0150833
R7249 VDD.n3661 VDD.n3646 0.0150833
R7250 VDD.n3707 VDD.n3693 0.0150833
R7251 VDD.n3786 VDD.n3771 0.0150833
R7252 VDD.n3832 VDD.n3828 0.0150833
R7253 VDD.n3957 VDD.n3956 0.0150833
R7254 VDD.n3960 VDD.n3959 0.0150833
R7255 VDD.n4001 VDD.n3986 0.0150833
R7256 VDD.n4024 VDD.n4009 0.0150833
R7257 VDD.n4032 VDD.n4031 0.0150833
R7258 VDD.n4083 VDD.n4081 0.0150833
R7259 VDD.n4160 VDD.n4156 0.0150833
R7260 VDD.n4251 VDD.n4250 0.0150833
R7261 VDD.n4307 VDD.n4303 0.0150833
R7262 VDD.n4481 VDD.n4480 0.0150833
R7263 VDD.n4549 VDD.n4548 0.0150833
R7264 VDD.n4912 VDD.n4906 0.0150833
R7265 VDD.n4968 VDD.n4967 0.0150833
R7266 VDD.n4991 VDD.n4990 0.0150833
R7267 VDD.n5051 VDD.n5050 0.0150833
R7268 VDD.n5085 VDD.n5073 0.0150833
R7269 VDD.n3042 VDD.n3041 0.013
R7270 VDD.n3486 VDD.n3471 0.013
R7271 VDD.n3556 VDD.n3537 0.013
R7272 VDD.n3595 VDD.n3580 0.013
R7273 VDD.n3791 VDD.n3790 0.013
R7274 VDD.n3806 VDD.n3791 0.013
R7275 VDD.n3809 VDD.n3807 0.013
R7276 VDD.n3884 VDD.n3879 0.013
R7277 VDD.n3916 VDD.n3901 0.013
R7278 VDD.n3955 VDD.n3940 0.013
R7279 VDD.n4120 VDD.n4119 0.013
R7280 VDD.n4180 VDD.n4177 0.013
R7281 VDD.n4197 VDD.n4196 0.013
R7282 VDD.n4315 VDD.n4314 0.013
R7283 VDD.n4405 VDD.n4404 0.013
R7284 VDD.n4462 VDD.n4458 0.013
R7285 VDD.n4714 VDD.n4713 0.013
R7286 VDD.n4737 VDD.n4736 0.013
R7287 VDD.n4837 VDD.n4836 0.013
R7288 VDD.n4882 VDD.n4881 0.013
R7289 VDD.n5142 VDD.n5141 0.013
R7290 VDD.n5143 VDD.n5142 0.013
R7291 VDD.n154 VDD.n142 0.0115132
R7292 VDD.n3073 VDD.n3072 0.0109167
R7293 VDD.n3104 VDD.n3103 0.0109167
R7294 VDD.n3135 VDD.n3134 0.0109167
R7295 VDD.n3166 VDD.n3165 0.0109167
R7296 VDD.n3197 VDD.n3196 0.0109167
R7297 VDD.n3228 VDD.n3227 0.0109167
R7298 VDD.n3259 VDD.n3258 0.0109167
R7299 VDD.n3290 VDD.n3289 0.0109167
R7300 VDD.n3321 VDD.n3320 0.0109167
R7301 VDD.n3352 VDD.n3351 0.0109167
R7302 VDD.n3383 VDD.n3382 0.0109167
R7303 VDD.n3488 VDD.n3487 0.0109167
R7304 VDD.n3493 VDD.n3492 0.0109167
R7305 VDD.n3621 VDD.n3620 0.0109167
R7306 VDD.n3644 VDD.n3641 0.0109167
R7307 VDD.n3663 VDD.n3662 0.0109167
R7308 VDD.n3727 VDD.n3713 0.0109167
R7309 VDD.n3748 VDD.n3747 0.0109167
R7310 VDD.n3766 VDD.n3751 0.0109167
R7311 VDD.n3834 VDD.n3833 0.0109167
R7312 VDD.n3973 VDD.n3960 0.0109167
R7313 VDD.n3978 VDD.n3974 0.0109167
R7314 VDD.n4003 VDD.n4002 0.0109167
R7315 VDD.n4046 VDD.n4033 0.0109167
R7316 VDD.n4118 VDD.n4105 0.0109167
R7317 VDD.n4162 VDD.n4161 0.0109167
R7318 VDD.n4177 VDD.n4176 0.0109167
R7319 VDD.n4269 VDD.n4268 0.0109167
R7320 VDD.n4309 VDD.n4308 0.0109167
R7321 VDD.n4328 VDD.n4315 0.0109167
R7322 VDD.n4336 VDD.n4335 0.0109167
R7323 VDD.n4464 VDD.n4463 0.0109167
R7324 VDD.n4562 VDD.n4561 0.0109167
R7325 VDD.n4627 VDD.n4612 0.0109167
R7326 VDD.n4629 VDD.n4628 0.0109167
R7327 VDD.n4657 VDD.n4656 0.0109167
R7328 VDD.n4718 VDD.n4716 0.0109167
R7329 VDD.n4796 VDD.n4795 0.0109167
R7330 VDD.n4879 VDD.n4878 0.0109167
R7331 VDD.n4963 VDD.n4962 0.0109167
R7332 VDD.n4967 VDD.n4966 0.0109167
R7333 VDD.n5047 VDD.n5046 0.0109167
R7334 VDD.n5123 VDD.n5122 0.0109167
R7335 VDD.n5129 VDD.n5128 0.0109167
R7336 VDD.n156 VDD.n155 0.00972509
R7337 VDD.n154 VDD.n153 0.00931057
R7338 VDD.n3450 VDD.n3449 0.00883333
R7339 VDD.n3512 VDD.n3494 0.00883333
R7340 VDD.n3575 VDD.n3560 0.00883333
R7341 VDD.n3577 VDD.n3576 0.00883333
R7342 VDD.n3646 VDD.n3645 0.00883333
R7343 VDD.n3826 VDD.n3812 0.00883333
R7344 VDD.n3894 VDD.n3889 0.00883333
R7345 VDD.n3934 VDD.n3919 0.00883333
R7346 VDD.n4009 VDD.n4008 0.00883333
R7347 VDD.n4136 VDD.n4123 0.00883333
R7348 VDD.n4139 VDD.n4137 0.00883333
R7349 VDD.n4201 VDD.n4198 0.00883333
R7350 VDD.n4267 VDD.n4254 0.00883333
R7351 VDD.n4408 VDD.n4407 0.00883333
R7352 VDD.n4423 VDD.n4422 0.00883333
R7353 VDD.n4485 VDD.n4481 0.00883333
R7354 VDD.n4503 VDD.n4502 0.00883333
R7355 VDD.n4504 VDD.n4503 0.00883333
R7356 VDD.n4794 VDD.n4790 0.00883333
R7357 VDD.n4811 VDD.n4810 0.00883333
R7358 VDD.n4878 VDD.n4877 0.00883333
R7359 VDD.n4946 VDD.n4945 0.00883333
R7360 VDD.n5048 VDD.n5047 0.00883333
R7361 VDD.n5121 VDD.n5120 0.00883333
R7362 VDD.n155 VDD.n138 0.00788007
R7363 VDD.n3077 VDD.n3076 0.00675
R7364 VDD.n3108 VDD.n3107 0.00675
R7365 VDD.n3139 VDD.n3138 0.00675
R7366 VDD.n3170 VDD.n3169 0.00675
R7367 VDD.n3201 VDD.n3200 0.00675
R7368 VDD.n3232 VDD.n3231 0.00675
R7369 VDD.n3263 VDD.n3262 0.00675
R7370 VDD.n3294 VDD.n3293 0.00675
R7371 VDD.n3325 VDD.n3324 0.00675
R7372 VDD.n3356 VDD.n3355 0.00675
R7373 VDD.n3387 VDD.n3386 0.00675
R7374 VDD.n3005 VDD.n3004 0.00675
R7375 VDD.n3406 VDD.n3405 0.00675
R7376 VDD.n3520 VDD.n3519 0.00675
R7377 VDD.n3667 VDD.n3664 0.00675
R7378 VDD.n3686 VDD.n3685 0.00675
R7379 VDD.n3746 VDD.n3731 0.00675
R7380 VDD.n3828 VDD.n3827 0.00675
R7381 VDD.n3851 VDD.n3850 0.00675
R7382 VDD.n3857 VDD.n3856 0.00675
R7383 VDD.n3984 VDD.n3981 0.00675
R7384 VDD.n4026 VDD.n4025 0.00675
R7385 VDD.n4052 VDD.n4050 0.00675
R7386 VDD.n4065 VDD.n4053 0.00675
R7387 VDD.n4099 VDD.n4086 0.00675
R7388 VDD.n4182 VDD.n4181 0.00675
R7389 VDD.n4254 VDD.n4253 0.00675
R7390 VDD.n4283 VDD.n4272 0.00675
R7391 VDD.n4288 VDD.n4284 0.00675
R7392 VDD.n4330 VDD.n4329 0.00675
R7393 VDD.n4335 VDD.n4334 0.00675
R7394 VDD.n4349 VDD.n4337 0.00675
R7395 VDD.n4421 VDD.n4408 0.00675
R7396 VDD.n4487 VDD.n4486 0.00675
R7397 VDD.n4583 VDD.n4582 0.00675
R7398 VDD.n4633 VDD.n4632 0.00675
R7399 VDD.n4650 VDD.n4635 0.00675
R7400 VDD.n4652 VDD.n4651 0.00675
R7401 VDD.n4658 VDD.n4657 0.00675
R7402 VDD.n4713 VDD.n4712 0.00675
R7403 VDD.n4790 VDD.n4789 0.00675
R7404 VDD.n4819 VDD.n4818 0.00675
R7405 VDD.n4944 VDD.n4943 0.00675
R7406 VDD.n4961 VDD.n4946 0.00675
R7407 VDD.n4986 VDD.n4985 0.00675
R7408 VDD.n5012 VDD.n5011 0.00675
R7409 VDD.n5028 VDD.n5027 0.00675
R7410 VDD.n5148 VDD.n5147 0.00675
R7411 VDD.n108 VDD.n105 0.00669723
R7412 VDD.n124 VDD.n123 0.00606809
R7413 VDD.n123 VDD.n122 0.00606809
R7414 VDD.n113 VDD.n112 0.0052619
R7415 VDD.n97 VDD.n96 0.00481034
R7416 VDD.n101 VDD.n100 0.00481034
R7417 VDD.n3430 VDD.n3429 0.00466667
R7418 VDD.n3558 VDD.n3557 0.00466667
R7419 VDD.n3669 VDD.n3668 0.00466667
R7420 VDD.n3849 VDD.n3835 0.00466667
R7421 VDD.n3900 VDD.n3897 0.00466667
R7422 VDD.n3986 VDD.n3985 0.00466667
R7423 VDD.n4105 VDD.n4104 0.00466667
R7424 VDD.n4154 VDD.n4142 0.00466667
R7425 VDD.n4196 VDD.n4195 0.00466667
R7426 VDD.n4217 VDD.n4215 0.00466667
R7427 VDD.n4221 VDD.n4218 0.00466667
R7428 VDD.n4236 VDD.n4233 0.00466667
R7429 VDD.n4438 VDD.n4426 0.00466667
R7430 VDD.n4442 VDD.n4440 0.00466667
R7431 VDD.n4479 VDD.n4478 0.00466667
R7432 VDD.n4508 VDD.n4505 0.00466667
R7433 VDD.n4548 VDD.n4547 0.00466667
R7434 VDD.n4565 VDD.n4562 0.00466667
R7435 VDD.n4612 VDD.n4611 0.00466667
R7436 VDD.n4754 VDD.n4753 0.00466667
R7437 VDD.n4788 VDD.n4787 0.00466667
R7438 VDD.n4817 VDD.n4813 0.00466667
R7439 VDD.n4838 VDD.n4837 0.00466667
R7440 VDD.n4847 VDD.n4846 0.00466667
R7441 VDD.n4859 VDD.n4858 0.00466667
R7442 VDD.n5068 VDD.n5067 0.00466667
R7443 VDD.n5102 VDD.n5101 0.00466667
R7444 VDD.n5106 VDD.n5104 0.00466667
R7445 VDD.n5127 VDD.n5123 0.00466667
R7446 VDD.n5270 VDD.n5269 0.00466667
R7447 VDD.n125 VDD.n124 0.00284423
R7448 VDD.n1794 VDD.n1661 0.00283209
R7449 VDD.n3059 VDD.n3058 0.00258333
R7450 VDD.n3090 VDD.n3089 0.00258333
R7451 VDD.n3121 VDD.n3120 0.00258333
R7452 VDD.n3152 VDD.n3151 0.00258333
R7453 VDD.n3183 VDD.n3182 0.00258333
R7454 VDD.n3214 VDD.n3213 0.00258333
R7455 VDD.n3245 VDD.n3244 0.00258333
R7456 VDD.n3276 VDD.n3275 0.00258333
R7457 VDD.n3307 VDD.n3306 0.00258333
R7458 VDD.n3338 VDD.n3337 0.00258333
R7459 VDD.n3369 VDD.n3368 0.00258333
R7460 VDD.n3425 VDD.n3424 0.00258333
R7461 VDD.n3514 VDD.n3513 0.00258333
R7462 VDD.n3596 VDD.n3595 0.00258333
R7463 VDD.n3601 VDD.n3600 0.00258333
R7464 VDD.n3691 VDD.n3687 0.00258333
R7465 VDD.n3729 VDD.n3728 0.00258333
R7466 VDD.n3767 VDD.n3766 0.00258333
R7467 VDD.n3935 VDD.n3934 0.00258333
R7468 VDD.n3940 VDD.n3939 0.00258333
R7469 VDD.n4007 VDD.n4004 0.00258333
R7470 VDD.n4031 VDD.n4030 0.00258333
R7471 VDD.n4080 VDD.n4068 0.00258333
R7472 VDD.n4100 VDD.n4099 0.00258333
R7473 VDD.n4156 VDD.n4155 0.00258333
R7474 VDD.n4237 VDD.n4236 0.00258333
R7475 VDD.n4294 VDD.n4291 0.00258333
R7476 VDD.n4313 VDD.n4312 0.00258333
R7477 VDD.n4355 VDD.n4353 0.00258333
R7478 VDD.n4368 VDD.n4356 0.00258333
R7479 VDD.n4385 VDD.n4384 0.00258333
R7480 VDD.n4401 VDD.n4389 0.00258333
R7481 VDD.n4402 VDD.n4401 0.00258333
R7482 VDD.n4458 VDD.n4457 0.00258333
R7483 VDD.n4558 VDD.n4557 0.00258333
R7484 VDD.n4589 VDD.n4586 0.00258333
R7485 VDD.n4604 VDD.n4600 0.00258333
R7486 VDD.n4610 VDD.n4609 0.00258333
R7487 VDD.n4673 VDD.n4659 0.00258333
R7488 VDD.n4679 VDD.n4677 0.00258333
R7489 VDD.n4694 VDD.n4693 0.00258333
R7490 VDD.n4733 VDD.n4732 0.00258333
R7491 VDD.n4751 VDD.n4737 0.00258333
R7492 VDD.n4902 VDD.n4901 0.00258333
R7493 VDD.n4903 VDD.n4902 0.00258333
R7494 VDD.n4919 VDD.n4918 0.00258333
R7495 VDD.n4938 VDD.n4921 0.00258333
R7496 VDD.n4984 VDD.n4969 0.00258333
R7497 VDD.n4992 VDD.n4991 0.00258333
R7498 VDD.n5007 VDD.n5006 0.00258333
R7499 VDD.n5067 VDD.n5066 0.00258333
R7500 VDD.n5086 VDD.n5085 0.00258333
R7501 VDD.n96 VDD.n95 0.00193678
R7502 VDD.n105 VDD.n101 0.00193678
R7503 VDD.n1796 VDD.n90 0.00149601
R7504 VDD.n125 VDD.n121 0.00106697
R7505 VDD.n1207 VDD.n1206 0.00100688
R7506 VDD.n892 VDD.n125 0.00100003
R7507 VDD.n901 VDD.n892 0.000567
R7508 VDD.n892 VDD.n133 0.000567
R7509 VDD.n892 VDD.n891 0.000567
R7510 VDD.n901 VDD.n900 0.000528434
R7511 VDD.n121 VDD.n120 0.000528434
R7512 VDD.n133 VDD.n132 0.000528434
R7513 VDD.n891 VDD.n890 0.000528434
R7514 VDD.n127 VDD.n126 0.000501607
R7515 VDD.n6791 VDD.n6790 0.000500267
R7516 VDD.n155 VDD.n154 0.00050023
R7517 VDD.n1661 VDD.n1660 0.000500078
R7518 VDD.n1794 VDD.n1793 0.000500038
R7519 VDD.n1795 VDD.n1794 0.00050001
R7520 VOUT.n746 VOUT.t156 27.6955
R7521 VOUT.n737 VOUT.t239 27.6955
R7522 VOUT.n737 VOUT.t163 27.6955
R7523 VOUT.n728 VOUT.t247 27.6955
R7524 VOUT.n728 VOUT.t238 27.6955
R7525 VOUT.n719 VOUT.t287 27.6955
R7526 VOUT.n719 VOUT.t188 27.6955
R7527 VOUT.n710 VOUT.t222 27.6955
R7528 VOUT.n710 VOUT.t323 27.6955
R7529 VOUT.n701 VOUT.t317 27.6955
R7530 VOUT.n701 VOUT.t204 27.6955
R7531 VOUT.n692 VOUT.t244 27.6955
R7532 VOUT.n692 VOUT.t293 27.6955
R7533 VOUT.n683 VOUT.t193 27.6955
R7534 VOUT.n683 VOUT.t240 27.6955
R7535 VOUT.n674 VOUT.t321 27.6955
R7536 VOUT.n674 VOUT.t271 27.6955
R7537 VOUT.n665 VOUT.t221 27.6955
R7538 VOUT.n665 VOUT.t338 27.6955
R7539 VOUT.n656 VOUT.t145 27.6955
R7540 VOUT.n656 VOUT.t237 27.6955
R7541 VOUT.n647 VOUT.t192 27.6955
R7542 VOUT.n647 VOUT.t292 27.6955
R7543 VOUT.n638 VOUT.t243 27.6955
R7544 VOUT.n638 VOUT.t251 27.6955
R7545 VOUT.n629 VOUT.t168 27.6955
R7546 VOUT.n629 VOUT.t322 27.6955
R7547 VOUT.n620 VOUT.t161 27.6955
R7548 VOUT.n620 VOUT.t316 27.6955
R7549 VOUT.n611 VOUT.t263 27.6955
R7550 VOUT.n611 VOUT.t216 27.6955
R7551 VOUT.n602 VOUT.t183 27.6955
R7552 VOUT.n602 VOUT.t284 27.6955
R7553 VOUT.n593 VOUT.t180 27.6955
R7554 VOUT.n593 VOUT.t334 27.6955
R7555 VOUT.n584 VOUT.t286 27.6955
R7556 VOUT.n584 VOUT.t235 27.6955
R7557 VOUT.n575 VOUT.t153 27.6955
R7558 VOUT.n575 VOUT.t306 27.6955
R7559 VOUT.n566 VOUT.t253 27.6955
R7560 VOUT.n934 VOUT.t170 27.6955
R7561 VOUT.n925 VOUT.t255 27.6955
R7562 VOUT.n925 VOUT.t179 27.6955
R7563 VOUT.n916 VOUT.t262 27.6955
R7564 VOUT.n916 VOUT.t254 27.6955
R7565 VOUT.n907 VOUT.t308 27.6955
R7566 VOUT.n907 VOUT.t198 27.6955
R7567 VOUT.n898 VOUT.t236 27.6955
R7568 VOUT.n898 VOUT.t337 27.6955
R7569 VOUT.n889 VOUT.t330 27.6955
R7570 VOUT.n889 VOUT.t213 27.6955
R7571 VOUT.n880 VOUT.t259 27.6955
R7572 VOUT.n880 VOUT.t311 27.6955
R7573 VOUT.n871 VOUT.t201 27.6955
R7574 VOUT.n871 VOUT.t256 27.6955
R7575 VOUT.n862 VOUT.t333 27.6955
R7576 VOUT.n862 VOUT.t285 27.6955
R7577 VOUT.n853 VOUT.t234 27.6955
R7578 VOUT.n853 VOUT.t155 27.6955
R7579 VOUT.n844 VOUT.t159 27.6955
R7580 VOUT.n844 VOUT.t252 27.6955
R7581 VOUT.n835 VOUT.t200 27.6955
R7582 VOUT.n835 VOUT.t309 27.6955
R7583 VOUT.n826 VOUT.t257 27.6955
R7584 VOUT.n826 VOUT.t267 27.6955
R7585 VOUT.n817 VOUT.t181 27.6955
R7586 VOUT.n817 VOUT.t336 27.6955
R7587 VOUT.n808 VOUT.t176 27.6955
R7588 VOUT.n808 VOUT.t329 27.6955
R7589 VOUT.n799 VOUT.t281 27.6955
R7590 VOUT.n799 VOUT.t230 27.6955
R7591 VOUT.n790 VOUT.t195 27.6955
R7592 VOUT.n790 VOUT.t302 27.6955
R7593 VOUT.n781 VOUT.t190 27.6955
R7594 VOUT.n781 VOUT.t149 27.6955
R7595 VOUT.n772 VOUT.t303 27.6955
R7596 VOUT.n772 VOUT.t248 27.6955
R7597 VOUT.n763 VOUT.t165 27.6955
R7598 VOUT.n763 VOUT.t319 27.6955
R7599 VOUT.n754 VOUT.t270 27.6955
R7600 VOUT.n1122 VOUT.t182 27.6955
R7601 VOUT.n1113 VOUT.t268 27.6955
R7602 VOUT.n1113 VOUT.t187 27.6955
R7603 VOUT.n1104 VOUT.t278 27.6955
R7604 VOUT.n1104 VOUT.t266 27.6955
R7605 VOUT.n1095 VOUT.t320 27.6955
R7606 VOUT.n1095 VOUT.t209 27.6955
R7607 VOUT.n1086 VOUT.t249 27.6955
R7608 VOUT.n1086 VOUT.t151 27.6955
R7609 VOUT.n1077 VOUT.t143 27.6955
R7610 VOUT.n1077 VOUT.t226 27.6955
R7611 VOUT.n1068 VOUT.t276 27.6955
R7612 VOUT.n1068 VOUT.t327 27.6955
R7613 VOUT.n1059 VOUT.t212 27.6955
R7614 VOUT.n1059 VOUT.t269 27.6955
R7615 VOUT.n1050 VOUT.t147 27.6955
R7616 VOUT.n1050 VOUT.t298 27.6955
R7617 VOUT.n1041 VOUT.t246 27.6955
R7618 VOUT.n1041 VOUT.t162 27.6955
R7619 VOUT.n1032 VOUT.t171 27.6955
R7620 VOUT.n1032 VOUT.t265 27.6955
R7621 VOUT.n1023 VOUT.t211 27.6955
R7622 VOUT.n1023 VOUT.t326 27.6955
R7623 VOUT.n1014 VOUT.t275 27.6955
R7624 VOUT.n1014 VOUT.t282 27.6955
R7625 VOUT.n1005 VOUT.t191 27.6955
R7626 VOUT.n1005 VOUT.t150 27.6955
R7627 VOUT.n996 VOUT.t185 27.6955
R7628 VOUT.n996 VOUT.t142 27.6955
R7629 VOUT.n987 VOUT.t291 27.6955
R7630 VOUT.n987 VOUT.t242 27.6955
R7631 VOUT.n978 VOUT.t203 27.6955
R7632 VOUT.n978 VOUT.t314 27.6955
R7633 VOUT.n969 VOUT.t197 27.6955
R7634 VOUT.n969 VOUT.t160 27.6955
R7635 VOUT.n960 VOUT.t315 27.6955
R7636 VOUT.n960 VOUT.t261 27.6955
R7637 VOUT.n951 VOUT.t178 27.6955
R7638 VOUT.n951 VOUT.t332 27.6955
R7639 VOUT.n942 VOUT.t283 27.6955
R7640 VOUT.n1310 VOUT.t335 27.6955
R7641 VOUT.n1301 VOUT.t219 27.6955
R7642 VOUT.n1301 VOUT.t144 27.6955
R7643 VOUT.n1292 VOUT.t227 27.6955
R7644 VOUT.n1292 VOUT.t218 27.6955
R7645 VOUT.n1283 VOUT.t264 27.6955
R7646 VOUT.n1283 VOUT.t169 27.6955
R7647 VOUT.n1274 VOUT.t207 27.6955
R7648 VOUT.n1274 VOUT.t301 27.6955
R7649 VOUT.n1265 VOUT.t289 27.6955
R7650 VOUT.n1265 VOUT.t189 27.6955
R7651 VOUT.n1256 VOUT.t224 27.6955
R7652 VOUT.n1256 VOUT.t273 27.6955
R7653 VOUT.n1247 VOUT.t175 27.6955
R7654 VOUT.n1247 VOUT.t220 27.6955
R7655 VOUT.n1238 VOUT.t294 27.6955
R7656 VOUT.n1238 VOUT.t245 27.6955
R7657 VOUT.n1229 VOUT.t206 27.6955
R7658 VOUT.n1229 VOUT.t318 27.6955
R7659 VOUT.n1220 VOUT.t325 27.6955
R7660 VOUT.n1220 VOUT.t217 27.6955
R7661 VOUT.n1211 VOUT.t173 27.6955
R7662 VOUT.n1211 VOUT.t272 27.6955
R7663 VOUT.n1202 VOUT.t223 27.6955
R7664 VOUT.n1202 VOUT.t229 27.6955
R7665 VOUT.n1193 VOUT.t148 27.6955
R7666 VOUT.n1193 VOUT.t300 27.6955
R7667 VOUT.n1184 VOUT.t139 27.6955
R7668 VOUT.n1184 VOUT.t288 27.6955
R7669 VOUT.n1175 VOUT.t241 27.6955
R7670 VOUT.n1175 VOUT.t202 27.6955
R7671 VOUT.n1166 VOUT.t164 27.6955
R7672 VOUT.n1166 VOUT.t258 27.6955
R7673 VOUT.n1157 VOUT.t157 27.6955
R7674 VOUT.n1157 VOUT.t312 27.6955
R7675 VOUT.n1148 VOUT.t260 27.6955
R7676 VOUT.n1148 VOUT.t214 27.6955
R7677 VOUT.n1139 VOUT.t331 27.6955
R7678 VOUT.n1139 VOUT.t280 27.6955
R7679 VOUT.n1130 VOUT.t231 27.6955
R7680 VOUT.n1498 VOUT.t199 27.6955
R7681 VOUT.n1489 VOUT.t297 27.6955
R7682 VOUT.n1489 VOUT.t208 27.6955
R7683 VOUT.n1480 VOUT.t307 27.6955
R7684 VOUT.n1480 VOUT.t296 27.6955
R7685 VOUT.n1471 VOUT.t146 27.6955
R7686 VOUT.n1471 VOUT.t228 27.6955
R7687 VOUT.n1462 VOUT.t279 27.6955
R7688 VOUT.n1462 VOUT.t177 27.6955
R7689 VOUT.n1453 VOUT.t167 27.6955
R7690 VOUT.n1453 VOUT.t250 27.6955
R7691 VOUT.n1444 VOUT.t305 27.6955
R7692 VOUT.n1444 VOUT.t154 27.6955
R7693 VOUT.n1435 VOUT.t233 27.6955
R7694 VOUT.n1435 VOUT.t299 27.6955
R7695 VOUT.n1426 VOUT.t172 27.6955
R7696 VOUT.n1426 VOUT.t328 27.6955
R7697 VOUT.n1417 VOUT.t277 27.6955
R7698 VOUT.n1417 VOUT.t186 27.6955
R7699 VOUT.n1408 VOUT.t194 27.6955
R7700 VOUT.n1408 VOUT.t295 27.6955
R7701 VOUT.n1399 VOUT.t232 27.6955
R7702 VOUT.n1399 VOUT.t152 27.6955
R7703 VOUT.n1390 VOUT.t304 27.6955
R7704 VOUT.n1390 VOUT.t310 27.6955
R7705 VOUT.n1381 VOUT.t210 27.6955
R7706 VOUT.n1381 VOUT.t174 27.6955
R7707 VOUT.n1372 VOUT.t205 27.6955
R7708 VOUT.n1372 VOUT.t166 27.6955
R7709 VOUT.n1363 VOUT.t324 27.6955
R7710 VOUT.n1363 VOUT.t274 27.6955
R7711 VOUT.n1354 VOUT.t225 27.6955
R7712 VOUT.n1354 VOUT.t140 27.6955
R7713 VOUT.n1345 VOUT.t215 27.6955
R7714 VOUT.n1345 VOUT.t184 27.6955
R7715 VOUT.n1336 VOUT.t141 27.6955
R7716 VOUT.n1336 VOUT.t290 27.6955
R7717 VOUT.n1327 VOUT.t196 27.6955
R7718 VOUT.n1327 VOUT.t158 27.6955
R7719 VOUT.n1318 VOUT.t313 27.6955
R7720 VOUT.n1689 VOUT.t501 27.6955
R7721 VOUT.n1680 VOUT.t406 27.6955
R7722 VOUT.n1680 VOUT.t132 27.6955
R7723 VOUT.n1671 VOUT.t503 27.6955
R7724 VOUT.n1671 VOUT.t478 27.6955
R7725 VOUT.n1662 VOUT.t79 27.6955
R7726 VOUT.n1662 VOUT.t19 27.6955
R7727 VOUT.n1653 VOUT.t377 27.6955
R7728 VOUT.n1653 VOUT.t64 27.6955
R7729 VOUT.n1644 VOUT.t371 27.6955
R7730 VOUT.n1644 VOUT.t466 27.6955
R7731 VOUT.n1635 VOUT.t126 27.6955
R7732 VOUT.n1635 VOUT.t491 27.6955
R7733 VOUT.n1626 VOUT.t104 27.6955
R7734 VOUT.n1626 VOUT.t418 27.6955
R7735 VOUT.n1617 VOUT.t116 27.6955
R7736 VOUT.n1617 VOUT.t506 27.6955
R7737 VOUT.n1608 VOUT.t423 27.6955
R7738 VOUT.n1608 VOUT.t117 27.6955
R7739 VOUT.n1599 VOUT.t134 27.6955
R7740 VOUT.n1599 VOUT.t17 27.6955
R7741 VOUT.n1590 VOUT.t513 27.6955
R7742 VOUT.n1590 VOUT.t63 27.6955
R7743 VOUT.n1581 VOUT.t127 27.6955
R7744 VOUT.n1581 VOUT.t57 27.6955
R7745 VOUT.n1572 VOUT.t430 27.6955
R7746 VOUT.n1572 VOUT.t512 27.6955
R7747 VOUT.n1563 VOUT.t21 27.6955
R7748 VOUT.n1563 VOUT.t374 27.6955
R7749 VOUT.n1554 VOUT.t389 27.6955
R7750 VOUT.n1554 VOUT.t42 27.6955
R7751 VOUT.n1545 VOUT.t52 27.6955
R7752 VOUT.n1545 VOUT.t355 27.6955
R7753 VOUT.n1536 VOUT.t393 27.6955
R7754 VOUT.n1536 VOUT.t490 27.6955
R7755 VOUT.n1527 VOUT.t78 27.6955
R7756 VOUT.n1527 VOUT.t397 27.6955
R7757 VOUT.n1518 VOUT.t369 27.6955
R7758 VOUT.n1518 VOUT.t357 27.6955
R7759 VOUT.n1509 VOUT.t45 27.6955
R7760 VOUT.n1874 VOUT.t440 27.6955
R7761 VOUT.n1865 VOUT.t487 27.6955
R7762 VOUT.n1865 VOUT.t34 27.6955
R7763 VOUT.n1856 VOUT.t120 27.6955
R7764 VOUT.n1856 VOUT.t366 27.6955
R7765 VOUT.n1847 VOUT.t489 27.6955
R7766 VOUT.n1847 VOUT.t427 27.6955
R7767 VOUT.n1838 VOUT.t118 27.6955
R7768 VOUT.n1838 VOUT.t68 27.6955
R7769 VOUT.n1829 VOUT.t5 27.6955
R7770 VOUT.n1829 VOUT.t29 27.6955
R7771 VOUT.n1820 VOUT.t114 27.6955
R7772 VOUT.n1820 VOUT.t73 27.6955
R7773 VOUT.n1811 VOUT.t13 27.6955
R7774 VOUT.n1811 VOUT.t388 27.6955
R7775 VOUT.n1802 VOUT.t40 27.6955
R7776 VOUT.n1802 VOUT.t497 27.6955
R7777 VOUT.n1793 VOUT.t342 27.6955
R7778 VOUT.n1793 VOUT.t27 27.6955
R7779 VOUT.n1784 VOUT.t351 27.6955
R7780 VOUT.n1784 VOUT.t23 27.6955
R7781 VOUT.n1775 VOUT.t414 27.6955
R7782 VOUT.n1775 VOUT.t500 27.6955
R7783 VOUT.n1766 VOUT.t24 27.6955
R7784 VOUT.n1766 VOUT.t61 27.6955
R7785 VOUT.n1757 VOUT.t441 27.6955
R7786 VOUT.n1757 VOUT.t375 27.6955
R7787 VOUT.n1748 VOUT.t75 27.6955
R7788 VOUT.n1748 VOUT.t379 27.6955
R7789 VOUT.n1739 VOUT.t76 27.6955
R7790 VOUT.n1739 VOUT.t88 27.6955
R7791 VOUT.n1730 VOUT.t412 27.6955
R7792 VOUT.n1730 VOUT.t59 27.6955
R7793 VOUT.n1721 VOUT.t404 27.6955
R7794 VOUT.n1721 VOUT.t66 27.6955
R7795 VOUT.n1712 VOUT.t130 27.6955
R7796 VOUT.n1712 VOUT.t62 27.6955
R7797 VOUT.n1703 VOUT.t422 27.6955
R7798 VOUT.n1703 VOUT.t105 27.6955
R7799 VOUT.n1694 VOUT.t22 27.6955
R7800 VOUT.n2062 VOUT.t385 27.6955
R7801 VOUT.n2053 VOUT.t494 27.6955
R7802 VOUT.n2053 VOUT.t386 27.6955
R7803 VOUT.n2044 VOUT.t37 27.6955
R7804 VOUT.n2044 VOUT.t109 27.6955
R7805 VOUT.n2035 VOUT.t25 27.6955
R7806 VOUT.n2035 VOUT.t349 27.6955
R7807 VOUT.n2026 VOUT.t391 27.6955
R7808 VOUT.n2026 VOUT.t384 27.6955
R7809 VOUT.n2017 VOUT.t46 27.6955
R7810 VOUT.n2017 VOUT.t51 27.6955
R7811 VOUT.n2008 VOUT.t438 27.6955
R7812 VOUT.n2008 VOUT.t92 27.6955
R7813 VOUT.n1999 VOUT.t103 27.6955
R7814 VOUT.n1999 VOUT.t350 27.6955
R7815 VOUT.n1990 VOUT.t47 27.6955
R7816 VOUT.n1990 VOUT.t492 27.6955
R7817 VOUT.n1981 VOUT.t421 27.6955
R7818 VOUT.n1981 VOUT.t96 27.6955
R7819 VOUT.n1972 VOUT.t121 27.6955
R7820 VOUT.n1972 VOUT.t413 27.6955
R7821 VOUT.n1963 VOUT.t106 27.6955
R7822 VOUT.n1963 VOUT.t81 27.6955
R7823 VOUT.n1954 VOUT.t394 27.6955
R7824 VOUT.n1954 VOUT.t464 27.6955
R7825 VOUT.n1945 VOUT.t100 27.6955
R7826 VOUT.n1945 VOUT.t48 27.6955
R7827 VOUT.n1936 VOUT.t122 27.6955
R7828 VOUT.n1936 VOUT.t94 27.6955
R7829 VOUT.n1927 VOUT.t93 27.6955
R7830 VOUT.n1927 VOUT.t483 27.6955
R7831 VOUT.n1918 VOUT.t91 27.6955
R7832 VOUT.n1918 VOUT.t390 27.6955
R7833 VOUT.n1909 VOUT.t368 27.6955
R7834 VOUT.n1909 VOUT.t131 27.6955
R7835 VOUT.n1900 VOUT.t361 27.6955
R7836 VOUT.n1900 VOUT.t415 27.6955
R7837 VOUT.n1891 VOUT.t95 27.6955
R7838 VOUT.n1891 VOUT.t488 27.6955
R7839 VOUT.n1882 VOUT.t87 27.6955
R7840 VOUT.n2250 VOUT.t425 27.6955
R7841 VOUT.n2241 VOUT.t44 27.6955
R7842 VOUT.n2241 VOUT.t381 27.6955
R7843 VOUT.n2232 VOUT.t82 27.6955
R7844 VOUT.n2232 VOUT.t71 27.6955
R7845 VOUT.n2223 VOUT.t376 27.6955
R7846 VOUT.n2223 VOUT.t340 27.6955
R7847 VOUT.n2214 VOUT.t123 27.6955
R7848 VOUT.n2214 VOUT.t101 27.6955
R7849 VOUT.n2205 VOUT.t462 27.6955
R7850 VOUT.n2205 VOUT.t3 27.6955
R7851 VOUT.n2196 VOUT.t498 27.6955
R7852 VOUT.n2196 VOUT.t133 27.6955
R7853 VOUT.n2187 VOUT.t395 27.6955
R7854 VOUT.n2187 VOUT.t486 27.6955
R7855 VOUT.n2178 VOUT.t463 27.6955
R7856 VOUT.n2178 VOUT.t124 27.6955
R7857 VOUT.n2169 VOUT.t110 27.6955
R7858 VOUT.n2169 VOUT.t56 27.6955
R7859 VOUT.n2160 VOUT.t85 27.6955
R7860 VOUT.n2160 VOUT.t119 27.6955
R7861 VOUT.n2151 VOUT.t129 27.6955
R7862 VOUT.n2151 VOUT.t67 27.6955
R7863 VOUT.n2142 VOUT.t72 27.6955
R7864 VOUT.n2142 VOUT.t370 27.6955
R7865 VOUT.n2133 VOUT.t90 27.6955
R7866 VOUT.n2133 VOUT.t41 27.6955
R7867 VOUT.n2124 VOUT.t429 27.6955
R7868 VOUT.n2124 VOUT.t353 27.6955
R7869 VOUT.n2115 VOUT.t74 27.6955
R7870 VOUT.n2115 VOUT.t356 27.6955
R7871 VOUT.n2106 VOUT.t428 27.6955
R7872 VOUT.n2106 VOUT.t499 27.6955
R7873 VOUT.n2097 VOUT.t419 27.6955
R7874 VOUT.n2097 VOUT.t485 27.6955
R7875 VOUT.n2088 VOUT.t502 27.6955
R7876 VOUT.n2088 VOUT.t372 27.6955
R7877 VOUT.n2079 VOUT.t102 27.6955
R7878 VOUT.n2079 VOUT.t493 27.6955
R7879 VOUT.n2070 VOUT.t26 27.6955
R7880 VOUT.n2258 VOUT.t8 27.6955
R7881 VOUT.n2265 VOUT.t496 27.6955
R7882 VOUT.n2265 VOUT.t32 27.6955
R7883 VOUT.n2272 VOUT.t80 27.6955
R7884 VOUT.n2272 VOUT.t505 27.6955
R7885 VOUT.n2279 VOUT.t507 27.6955
R7886 VOUT.n2279 VOUT.t363 27.6955
R7887 VOUT.n2286 VOUT.t125 27.6955
R7888 VOUT.n2286 VOUT.t378 27.6955
R7889 VOUT.n2293 VOUT.t65 27.6955
R7890 VOUT.n2293 VOUT.t12 27.6955
R7891 VOUT.n2300 VOUT.t20 27.6955
R7892 VOUT.n2300 VOUT.t112 27.6955
R7893 VOUT.n2307 VOUT.t70 27.6955
R7894 VOUT.n2307 VOUT.t58 27.6955
R7895 VOUT.n2314 VOUT.t39 27.6955
R7896 VOUT.n2314 VOUT.t111 27.6955
R7897 VOUT.n2321 VOUT.t352 27.6955
R7898 VOUT.n2321 VOUT.t509 27.6955
R7899 VOUT.n2328 VOUT.t508 27.6955
R7900 VOUT.n2328 VOUT.t373 27.6955
R7901 VOUT.n2335 VOUT.t107 27.6955
R7902 VOUT.n2335 VOUT.t99 27.6955
R7903 VOUT.n2342 VOUT.t364 27.6955
R7904 VOUT.n2342 VOUT.t77 27.6955
R7905 VOUT.n2349 VOUT.t343 27.6955
R7906 VOUT.n2349 VOUT.t344 27.6955
R7907 VOUT.n2356 VOUT.t86 27.6955
R7908 VOUT.n2356 VOUT.t367 27.6955
R7909 VOUT.n2363 VOUT.t495 27.6955
R7910 VOUT.n2363 VOUT.t18 27.6955
R7911 VOUT.n2370 VOUT.t9 27.6955
R7912 VOUT.n2370 VOUT.t4 27.6955
R7913 VOUT.n2377 VOUT.t405 27.6955
R7914 VOUT.n2377 VOUT.t83 27.6955
R7915 VOUT.n2384 VOUT.t115 27.6955
R7916 VOUT.n2384 VOUT.t504 27.6955
R7917 VOUT.n2391 VOUT.t358 27.6955
R7918 VOUT.n2391 VOUT.t98 27.6955
R7919 VOUT.n2398 VOUT.t365 27.6955
R7920 VOUT.n556 VOUT.t460 16.5305
R7921 VOUT.n547 VOUT.t468 16.5305
R7922 VOUT.n547 VOUT.t411 16.5305
R7923 VOUT.n538 VOUT.t453 16.5305
R7924 VOUT.n538 VOUT.t1 16.5305
R7925 VOUT.n529 VOUT.t113 16.5305
R7926 VOUT.n529 VOUT.t400 16.5305
R7927 VOUT.n520 VOUT.t469 16.5305
R7928 VOUT.n520 VOUT.t482 16.5305
R7929 VOUT.n511 VOUT.t7 16.5305
R7930 VOUT.n511 VOUT.t399 16.5305
R7931 VOUT.n502 VOUT.t16 16.5305
R7932 VOUT.n502 VOUT.t519 16.5305
R7933 VOUT.n493 VOUT.t392 16.5305
R7934 VOUT.n493 VOUT.t437 16.5305
R7935 VOUT.n484 VOUT.t511 16.5305
R7936 VOUT.n484 VOUT.t471 16.5305
R7937 VOUT.n475 VOUT.t446 16.5305
R7938 VOUT.n475 VOUT.t138 16.5305
R7939 VOUT.n466 VOUT.t442 16.5305
R7940 VOUT.n466 VOUT.t6 16.5305
R7941 VOUT.n457 VOUT.t455 16.5305
R7942 VOUT.n457 VOUT.t348 16.5305
R7943 VOUT.n448 VOUT.t474 16.5305
R7944 VOUT.n448 VOUT.t401 16.5305
R7945 VOUT.n439 VOUT.t450 16.5305
R7946 VOUT.n439 VOUT.t15 16.5305
R7947 VOUT.n430 VOUT.t345 16.5305
R7948 VOUT.n430 VOUT.t458 16.5305
R7949 VOUT.n421 VOUT.t55 16.5305
R7950 VOUT.n421 VOUT.t439 16.5305
R7951 VOUT.n412 VOUT.t467 16.5305
R7952 VOUT.n412 VOUT.t11 16.5305
R7953 VOUT.n403 VOUT.t360 16.5305
R7954 VOUT.n403 VOUT.t38 16.5305
R7955 VOUT.n394 VOUT.t476 16.5305
R7956 VOUT.n394 VOUT.t398 16.5305
R7957 VOUT.n385 VOUT.t470 16.5305
R7958 VOUT.n385 VOUT.t461 16.5305
R7959 VOUT.n377 VOUT.t475 16.5305
R7960 VOUT.n368 VOUT.t518 16.5305
R7961 VOUT.n359 VOUT.t403 16.5305
R7962 VOUT.n359 VOUT.t43 16.5305
R7963 VOUT.n350 VOUT.t443 16.5305
R7964 VOUT.n350 VOUT.t135 16.5305
R7965 VOUT.n341 VOUT.t409 16.5305
R7966 VOUT.n341 VOUT.t416 16.5305
R7967 VOUT.n332 VOUT.t480 16.5305
R7968 VOUT.n332 VOUT.t137 16.5305
R7969 VOUT.n323 VOUT.t33 16.5305
R7970 VOUT.n323 VOUT.t54 16.5305
R7971 VOUT.n314 VOUT.t516 16.5305
R7972 VOUT.n314 VOUT.t408 16.5305
R7973 VOUT.n305 VOUT.t69 16.5305
R7974 VOUT.n305 VOUT.t346 16.5305
R7975 VOUT.n296 VOUT.t36 16.5305
R7976 VOUT.n296 VOUT.t432 16.5305
R7977 VOUT.n287 VOUT.t515 16.5305
R7978 VOUT.n287 VOUT.t60 16.5305
R7979 VOUT.n278 VOUT.t128 16.5305
R7980 VOUT.n278 VOUT.t28 16.5305
R7981 VOUT.n269 VOUT.t457 16.5305
R7982 VOUT.n269 VOUT.t420 16.5305
R7983 VOUT.n260 VOUT.t359 16.5305
R7984 VOUT.n260 VOUT.t433 16.5305
R7985 VOUT.n251 VOUT.t434 16.5305
R7986 VOUT.n251 VOUT.t380 16.5305
R7987 VOUT.n242 VOUT.t417 16.5305
R7988 VOUT.n242 VOUT.t445 16.5305
R7989 VOUT.n233 VOUT.t517 16.5305
R7990 VOUT.n233 VOUT.t341 16.5305
R7991 VOUT.n224 VOUT.t339 16.5305
R7992 VOUT.n224 VOUT.t436 16.5305
R7993 VOUT.n215 VOUT.t396 16.5305
R7994 VOUT.n215 VOUT.t97 16.5305
R7995 VOUT.n206 VOUT.t456 16.5305
R7996 VOUT.n206 VOUT.t14 16.5305
R7997 VOUT.n197 VOUT.t510 16.5305
R7998 VOUT.n197 VOUT.t454 16.5305
R7999 VOUT.n189 VOUT.t451 16.5305
R8000 VOUT.n180 VOUT.t49 16.5305
R8001 VOUT.n171 VOUT.t347 16.5305
R8002 VOUT.n171 VOUT.t449 16.5305
R8003 VOUT.n162 VOUT.t30 16.5305
R8004 VOUT.n162 VOUT.t424 16.5305
R8005 VOUT.n153 VOUT.t0 16.5305
R8006 VOUT.n153 VOUT.t136 16.5305
R8007 VOUT.n144 VOUT.t410 16.5305
R8008 VOUT.n144 VOUT.t473 16.5305
R8009 VOUT.n135 VOUT.t108 16.5305
R8010 VOUT.n135 VOUT.t383 16.5305
R8011 VOUT.n126 VOUT.t382 16.5305
R8012 VOUT.n126 VOUT.t402 16.5305
R8013 VOUT.n117 VOUT.t10 16.5305
R8014 VOUT.n117 VOUT.t2 16.5305
R8015 VOUT.n108 VOUT.t477 16.5305
R8016 VOUT.n108 VOUT.t484 16.5305
R8017 VOUT.n99 VOUT.t426 16.5305
R8018 VOUT.n99 VOUT.t407 16.5305
R8019 VOUT.n90 VOUT.t444 16.5305
R8020 VOUT.n90 VOUT.t50 16.5305
R8021 VOUT.n81 VOUT.t89 16.5305
R8022 VOUT.n81 VOUT.t35 16.5305
R8023 VOUT.n72 VOUT.t435 16.5305
R8024 VOUT.n72 VOUT.t31 16.5305
R8025 VOUT.n63 VOUT.t479 16.5305
R8026 VOUT.n63 VOUT.t447 16.5305
R8027 VOUT.n54 VOUT.t84 16.5305
R8028 VOUT.n54 VOUT.t354 16.5305
R8029 VOUT.n45 VOUT.t448 16.5305
R8030 VOUT.n45 VOUT.t452 16.5305
R8031 VOUT.n36 VOUT.t53 16.5305
R8032 VOUT.n36 VOUT.t431 16.5305
R8033 VOUT.n27 VOUT.t459 16.5305
R8034 VOUT.n27 VOUT.t387 16.5305
R8035 VOUT.n18 VOUT.t362 16.5305
R8036 VOUT.n18 VOUT.t472 16.5305
R8037 VOUT.n9 VOUT.t514 16.5305
R8038 VOUT.n9 VOUT.t465 16.5305
R8039 VOUT.n1 VOUT.t481 16.5305
R8040 VOUT.n2259 VOUT.n2258 13.1521
R8041 VOUT.n2399 VOUT.n2398 13.1521
R8042 VOUT.n2266 VOUT.n2265 13.1512
R8043 VOUT.n2273 VOUT.n2272 13.1512
R8044 VOUT.n2280 VOUT.n2279 13.1512
R8045 VOUT.n2287 VOUT.n2286 13.1512
R8046 VOUT.n2294 VOUT.n2293 13.1512
R8047 VOUT.n2301 VOUT.n2300 13.1512
R8048 VOUT.n2308 VOUT.n2307 13.1512
R8049 VOUT.n2315 VOUT.n2314 13.1512
R8050 VOUT.n2322 VOUT.n2321 13.1512
R8051 VOUT.n2329 VOUT.n2328 13.1512
R8052 VOUT.n2336 VOUT.n2335 13.1512
R8053 VOUT.n2343 VOUT.n2342 13.1512
R8054 VOUT.n2350 VOUT.n2349 13.1512
R8055 VOUT.n2357 VOUT.n2356 13.1512
R8056 VOUT.n2364 VOUT.n2363 13.1512
R8057 VOUT.n2371 VOUT.n2370 13.1512
R8058 VOUT.n2378 VOUT.n2377 13.1512
R8059 VOUT.n2385 VOUT.n2384 13.1512
R8060 VOUT.n2392 VOUT.n2391 13.1512
R8061 VOUT.n2251 VOUT.n2250 13.149
R8062 VOUT.n2071 VOUT.n2070 13.149
R8063 VOUT.n2242 VOUT.n2241 13.1481
R8064 VOUT.n2233 VOUT.n2232 13.1481
R8065 VOUT.n2224 VOUT.n2223 13.1481
R8066 VOUT.n2215 VOUT.n2214 13.1481
R8067 VOUT.n2206 VOUT.n2205 13.1481
R8068 VOUT.n2197 VOUT.n2196 13.1481
R8069 VOUT.n2188 VOUT.n2187 13.1481
R8070 VOUT.n2179 VOUT.n2178 13.1481
R8071 VOUT.n2170 VOUT.n2169 13.1481
R8072 VOUT.n2161 VOUT.n2160 13.1481
R8073 VOUT.n2152 VOUT.n2151 13.1481
R8074 VOUT.n2143 VOUT.n2142 13.1481
R8075 VOUT.n2134 VOUT.n2133 13.1481
R8076 VOUT.n2125 VOUT.n2124 13.1481
R8077 VOUT.n2116 VOUT.n2115 13.1481
R8078 VOUT.n2107 VOUT.n2106 13.1481
R8079 VOUT.n2098 VOUT.n2097 13.1481
R8080 VOUT.n2089 VOUT.n2088 13.1481
R8081 VOUT.n2080 VOUT.n2079 13.1481
R8082 VOUT.n1875 VOUT.n1874 13.1451
R8083 VOUT.n1695 VOUT.n1694 13.1451
R8084 VOUT.n1866 VOUT.n1865 13.1442
R8085 VOUT.n1857 VOUT.n1856 13.1442
R8086 VOUT.n1848 VOUT.n1847 13.1442
R8087 VOUT.n1839 VOUT.n1838 13.1442
R8088 VOUT.n1830 VOUT.n1829 13.1442
R8089 VOUT.n1821 VOUT.n1820 13.1442
R8090 VOUT.n1812 VOUT.n1811 13.1442
R8091 VOUT.n1803 VOUT.n1802 13.1442
R8092 VOUT.n1794 VOUT.n1793 13.1442
R8093 VOUT.n1785 VOUT.n1784 13.1442
R8094 VOUT.n1776 VOUT.n1775 13.1442
R8095 VOUT.n1767 VOUT.n1766 13.1442
R8096 VOUT.n1758 VOUT.n1757 13.1442
R8097 VOUT.n1749 VOUT.n1748 13.1442
R8098 VOUT.n1740 VOUT.n1739 13.1442
R8099 VOUT.n1731 VOUT.n1730 13.1442
R8100 VOUT.n1722 VOUT.n1721 13.1442
R8101 VOUT.n1713 VOUT.n1712 13.1442
R8102 VOUT.n1704 VOUT.n1703 13.1442
R8103 VOUT.n747 VOUT.n746 13.1434
R8104 VOUT.n567 VOUT.n566 13.1434
R8105 VOUT.n2063 VOUT.n2062 13.1434
R8106 VOUT.n1883 VOUT.n1882 13.1434
R8107 VOUT.n738 VOUT.n737 13.1425
R8108 VOUT.n729 VOUT.n728 13.1425
R8109 VOUT.n720 VOUT.n719 13.1425
R8110 VOUT.n711 VOUT.n710 13.1425
R8111 VOUT.n702 VOUT.n701 13.1425
R8112 VOUT.n693 VOUT.n692 13.1425
R8113 VOUT.n684 VOUT.n683 13.1425
R8114 VOUT.n675 VOUT.n674 13.1425
R8115 VOUT.n666 VOUT.n665 13.1425
R8116 VOUT.n657 VOUT.n656 13.1425
R8117 VOUT.n648 VOUT.n647 13.1425
R8118 VOUT.n639 VOUT.n638 13.1425
R8119 VOUT.n630 VOUT.n629 13.1425
R8120 VOUT.n621 VOUT.n620 13.1425
R8121 VOUT.n612 VOUT.n611 13.1425
R8122 VOUT.n603 VOUT.n602 13.1425
R8123 VOUT.n594 VOUT.n593 13.1425
R8124 VOUT.n585 VOUT.n584 13.1425
R8125 VOUT.n576 VOUT.n575 13.1425
R8126 VOUT.n2054 VOUT.n2053 13.1425
R8127 VOUT.n2045 VOUT.n2044 13.1425
R8128 VOUT.n2036 VOUT.n2035 13.1425
R8129 VOUT.n2027 VOUT.n2026 13.1425
R8130 VOUT.n2018 VOUT.n2017 13.1425
R8131 VOUT.n2009 VOUT.n2008 13.1425
R8132 VOUT.n2000 VOUT.n1999 13.1425
R8133 VOUT.n1991 VOUT.n1990 13.1425
R8134 VOUT.n1982 VOUT.n1981 13.1425
R8135 VOUT.n1973 VOUT.n1972 13.1425
R8136 VOUT.n1964 VOUT.n1963 13.1425
R8137 VOUT.n1955 VOUT.n1954 13.1425
R8138 VOUT.n1946 VOUT.n1945 13.1425
R8139 VOUT.n1937 VOUT.n1936 13.1425
R8140 VOUT.n1928 VOUT.n1927 13.1425
R8141 VOUT.n1919 VOUT.n1918 13.1425
R8142 VOUT.n1910 VOUT.n1909 13.1425
R8143 VOUT.n1901 VOUT.n1900 13.1425
R8144 VOUT.n1892 VOUT.n1891 13.1425
R8145 VOUT.n935 VOUT.n934 13.1422
R8146 VOUT.n755 VOUT.n754 13.1422
R8147 VOUT.n926 VOUT.n925 13.1413
R8148 VOUT.n917 VOUT.n916 13.1413
R8149 VOUT.n908 VOUT.n907 13.1413
R8150 VOUT.n899 VOUT.n898 13.1413
R8151 VOUT.n890 VOUT.n889 13.1413
R8152 VOUT.n881 VOUT.n880 13.1413
R8153 VOUT.n872 VOUT.n871 13.1413
R8154 VOUT.n863 VOUT.n862 13.1413
R8155 VOUT.n854 VOUT.n853 13.1413
R8156 VOUT.n845 VOUT.n844 13.1413
R8157 VOUT.n836 VOUT.n835 13.1413
R8158 VOUT.n827 VOUT.n826 13.1413
R8159 VOUT.n818 VOUT.n817 13.1413
R8160 VOUT.n809 VOUT.n808 13.1413
R8161 VOUT.n800 VOUT.n799 13.1413
R8162 VOUT.n791 VOUT.n790 13.1413
R8163 VOUT.n782 VOUT.n781 13.1413
R8164 VOUT.n773 VOUT.n772 13.1413
R8165 VOUT.n764 VOUT.n763 13.1413
R8166 VOUT.n1123 VOUT.n1122 13.1402
R8167 VOUT.n943 VOUT.n942 13.1402
R8168 VOUT.n1114 VOUT.n1113 13.1393
R8169 VOUT.n1105 VOUT.n1104 13.1393
R8170 VOUT.n1096 VOUT.n1095 13.1393
R8171 VOUT.n1087 VOUT.n1086 13.1393
R8172 VOUT.n1078 VOUT.n1077 13.1393
R8173 VOUT.n1069 VOUT.n1068 13.1393
R8174 VOUT.n1060 VOUT.n1059 13.1393
R8175 VOUT.n1051 VOUT.n1050 13.1393
R8176 VOUT.n1042 VOUT.n1041 13.1393
R8177 VOUT.n1033 VOUT.n1032 13.1393
R8178 VOUT.n1024 VOUT.n1023 13.1393
R8179 VOUT.n1015 VOUT.n1014 13.1393
R8180 VOUT.n1006 VOUT.n1005 13.1393
R8181 VOUT.n997 VOUT.n996 13.1393
R8182 VOUT.n988 VOUT.n987 13.1393
R8183 VOUT.n979 VOUT.n978 13.1393
R8184 VOUT.n970 VOUT.n969 13.1393
R8185 VOUT.n961 VOUT.n960 13.1393
R8186 VOUT.n952 VOUT.n951 13.1393
R8187 VOUT.n1311 VOUT.n1310 13.1381
R8188 VOUT.n1131 VOUT.n1130 13.1381
R8189 VOUT.n1302 VOUT.n1301 13.1372
R8190 VOUT.n1293 VOUT.n1292 13.1372
R8191 VOUT.n1284 VOUT.n1283 13.1372
R8192 VOUT.n1275 VOUT.n1274 13.1372
R8193 VOUT.n1266 VOUT.n1265 13.1372
R8194 VOUT.n1257 VOUT.n1256 13.1372
R8195 VOUT.n1248 VOUT.n1247 13.1372
R8196 VOUT.n1239 VOUT.n1238 13.1372
R8197 VOUT.n1230 VOUT.n1229 13.1372
R8198 VOUT.n1221 VOUT.n1220 13.1372
R8199 VOUT.n1212 VOUT.n1211 13.1372
R8200 VOUT.n1203 VOUT.n1202 13.1372
R8201 VOUT.n1194 VOUT.n1193 13.1372
R8202 VOUT.n1185 VOUT.n1184 13.1372
R8203 VOUT.n1176 VOUT.n1175 13.1372
R8204 VOUT.n1167 VOUT.n1166 13.1372
R8205 VOUT.n1158 VOUT.n1157 13.1372
R8206 VOUT.n1149 VOUT.n1148 13.1372
R8207 VOUT.n1140 VOUT.n1139 13.1372
R8208 VOUT.n1499 VOUT.n1498 13.1359
R8209 VOUT.n1319 VOUT.n1318 13.1359
R8210 VOUT.n1490 VOUT.n1489 13.135
R8211 VOUT.n1481 VOUT.n1480 13.135
R8212 VOUT.n1472 VOUT.n1471 13.135
R8213 VOUT.n1463 VOUT.n1462 13.135
R8214 VOUT.n1454 VOUT.n1453 13.135
R8215 VOUT.n1445 VOUT.n1444 13.135
R8216 VOUT.n1436 VOUT.n1435 13.135
R8217 VOUT.n1427 VOUT.n1426 13.135
R8218 VOUT.n1418 VOUT.n1417 13.135
R8219 VOUT.n1409 VOUT.n1408 13.135
R8220 VOUT.n1400 VOUT.n1399 13.135
R8221 VOUT.n1391 VOUT.n1390 13.135
R8222 VOUT.n1382 VOUT.n1381 13.135
R8223 VOUT.n1373 VOUT.n1372 13.135
R8224 VOUT.n1364 VOUT.n1363 13.135
R8225 VOUT.n1355 VOUT.n1354 13.135
R8226 VOUT.n1346 VOUT.n1345 13.135
R8227 VOUT.n1337 VOUT.n1336 13.135
R8228 VOUT.n1328 VOUT.n1327 13.135
R8229 VOUT.n557 VOUT.n556 11.6601
R8230 VOUT.n548 VOUT.n547 11.6601
R8231 VOUT.n539 VOUT.n538 11.6601
R8232 VOUT.n530 VOUT.n529 11.6601
R8233 VOUT.n521 VOUT.n520 11.6601
R8234 VOUT.n512 VOUT.n511 11.6601
R8235 VOUT.n503 VOUT.n502 11.6601
R8236 VOUT.n494 VOUT.n493 11.6601
R8237 VOUT.n485 VOUT.n484 11.6601
R8238 VOUT.n476 VOUT.n475 11.6601
R8239 VOUT.n467 VOUT.n466 11.6601
R8240 VOUT.n458 VOUT.n457 11.6601
R8241 VOUT.n449 VOUT.n448 11.6601
R8242 VOUT.n440 VOUT.n439 11.6601
R8243 VOUT.n431 VOUT.n430 11.6601
R8244 VOUT.n422 VOUT.n421 11.6601
R8245 VOUT.n413 VOUT.n412 11.6601
R8246 VOUT.n404 VOUT.n403 11.6601
R8247 VOUT.n395 VOUT.n394 11.6601
R8248 VOUT.n386 VOUT.n385 11.6601
R8249 VOUT.n378 VOUT.n377 11.6601
R8250 VOUT.n369 VOUT.n368 11.6601
R8251 VOUT.n360 VOUT.n359 11.6601
R8252 VOUT.n351 VOUT.n350 11.6601
R8253 VOUT.n342 VOUT.n341 11.6601
R8254 VOUT.n333 VOUT.n332 11.6601
R8255 VOUT.n324 VOUT.n323 11.6601
R8256 VOUT.n315 VOUT.n314 11.6601
R8257 VOUT.n306 VOUT.n305 11.6601
R8258 VOUT.n297 VOUT.n296 11.6601
R8259 VOUT.n288 VOUT.n287 11.6601
R8260 VOUT.n279 VOUT.n278 11.6601
R8261 VOUT.n270 VOUT.n269 11.6601
R8262 VOUT.n261 VOUT.n260 11.6601
R8263 VOUT.n252 VOUT.n251 11.6601
R8264 VOUT.n243 VOUT.n242 11.6601
R8265 VOUT.n234 VOUT.n233 11.6601
R8266 VOUT.n225 VOUT.n224 11.6601
R8267 VOUT.n216 VOUT.n215 11.6601
R8268 VOUT.n207 VOUT.n206 11.6601
R8269 VOUT.n198 VOUT.n197 11.6601
R8270 VOUT.n190 VOUT.n189 11.6601
R8271 VOUT.n181 VOUT.n180 11.6601
R8272 VOUT.n172 VOUT.n171 11.6601
R8273 VOUT.n163 VOUT.n162 11.6601
R8274 VOUT.n154 VOUT.n153 11.6601
R8275 VOUT.n145 VOUT.n144 11.6601
R8276 VOUT.n136 VOUT.n135 11.6601
R8277 VOUT.n127 VOUT.n126 11.6601
R8278 VOUT.n118 VOUT.n117 11.6601
R8279 VOUT.n109 VOUT.n108 11.6601
R8280 VOUT.n100 VOUT.n99 11.6601
R8281 VOUT.n91 VOUT.n90 11.6601
R8282 VOUT.n82 VOUT.n81 11.6601
R8283 VOUT.n73 VOUT.n72 11.6601
R8284 VOUT.n64 VOUT.n63 11.6601
R8285 VOUT.n55 VOUT.n54 11.6601
R8286 VOUT.n46 VOUT.n45 11.6601
R8287 VOUT.n37 VOUT.n36 11.6601
R8288 VOUT.n28 VOUT.n27 11.6601
R8289 VOUT.n19 VOUT.n18 11.6601
R8290 VOUT.n10 VOUT.n9 11.6601
R8291 VOUT.n2 VOUT.n1 11.6601
R8292 VOUT.n1690 VOUT.n1689 9.02061
R8293 VOUT.n1681 VOUT.n1680 9.02061
R8294 VOUT.n1672 VOUT.n1671 9.02061
R8295 VOUT.n1663 VOUT.n1662 9.02061
R8296 VOUT.n1654 VOUT.n1653 9.02061
R8297 VOUT.n1645 VOUT.n1644 9.02061
R8298 VOUT.n1636 VOUT.n1635 9.02061
R8299 VOUT.n1627 VOUT.n1626 9.02061
R8300 VOUT.n1618 VOUT.n1617 9.02061
R8301 VOUT.n1609 VOUT.n1608 9.02061
R8302 VOUT.n1600 VOUT.n1599 9.02061
R8303 VOUT.n1591 VOUT.n1590 9.02061
R8304 VOUT.n1582 VOUT.n1581 9.02061
R8305 VOUT.n1573 VOUT.n1572 9.02061
R8306 VOUT.n1564 VOUT.n1563 9.02061
R8307 VOUT.n1555 VOUT.n1554 9.02061
R8308 VOUT.n1546 VOUT.n1545 9.02061
R8309 VOUT.n1537 VOUT.n1536 9.02061
R8310 VOUT.n1528 VOUT.n1527 9.02061
R8311 VOUT.n1519 VOUT.n1518 9.02061
R8312 VOUT.n1510 VOUT.n1509 9.02061
R8313 VOUT.n382 VOUT.n381 4.5005
R8314 VOUT.n390 VOUT.n389 4.5005
R8315 VOUT.n399 VOUT.n398 4.5005
R8316 VOUT.n408 VOUT.n407 4.5005
R8317 VOUT.n417 VOUT.n416 4.5005
R8318 VOUT.n426 VOUT.n425 4.5005
R8319 VOUT.n435 VOUT.n434 4.5005
R8320 VOUT.n444 VOUT.n443 4.5005
R8321 VOUT.n453 VOUT.n452 4.5005
R8322 VOUT.n462 VOUT.n461 4.5005
R8323 VOUT.n471 VOUT.n470 4.5005
R8324 VOUT.n480 VOUT.n479 4.5005
R8325 VOUT.n489 VOUT.n488 4.5005
R8326 VOUT.n498 VOUT.n497 4.5005
R8327 VOUT.n507 VOUT.n506 4.5005
R8328 VOUT.n516 VOUT.n515 4.5005
R8329 VOUT.n525 VOUT.n524 4.5005
R8330 VOUT.n534 VOUT.n533 4.5005
R8331 VOUT.n543 VOUT.n542 4.5005
R8332 VOUT.n552 VOUT.n551 4.5005
R8333 VOUT.n561 VOUT.n560 4.5005
R8334 VOUT.n194 VOUT.n193 4.5005
R8335 VOUT.n202 VOUT.n201 4.5005
R8336 VOUT.n211 VOUT.n210 4.5005
R8337 VOUT.n220 VOUT.n219 4.5005
R8338 VOUT.n229 VOUT.n228 4.5005
R8339 VOUT.n238 VOUT.n237 4.5005
R8340 VOUT.n247 VOUT.n246 4.5005
R8341 VOUT.n256 VOUT.n255 4.5005
R8342 VOUT.n265 VOUT.n264 4.5005
R8343 VOUT.n274 VOUT.n273 4.5005
R8344 VOUT.n283 VOUT.n282 4.5005
R8345 VOUT.n292 VOUT.n291 4.5005
R8346 VOUT.n301 VOUT.n300 4.5005
R8347 VOUT.n310 VOUT.n309 4.5005
R8348 VOUT.n319 VOUT.n318 4.5005
R8349 VOUT.n328 VOUT.n327 4.5005
R8350 VOUT.n337 VOUT.n336 4.5005
R8351 VOUT.n346 VOUT.n345 4.5005
R8352 VOUT.n355 VOUT.n354 4.5005
R8353 VOUT.n364 VOUT.n363 4.5005
R8354 VOUT.n373 VOUT.n372 4.5005
R8355 VOUT.n6 VOUT.n5 4.5005
R8356 VOUT.n14 VOUT.n13 4.5005
R8357 VOUT.n23 VOUT.n22 4.5005
R8358 VOUT.n32 VOUT.n31 4.5005
R8359 VOUT.n41 VOUT.n40 4.5005
R8360 VOUT.n50 VOUT.n49 4.5005
R8361 VOUT.n59 VOUT.n58 4.5005
R8362 VOUT.n68 VOUT.n67 4.5005
R8363 VOUT.n77 VOUT.n76 4.5005
R8364 VOUT.n86 VOUT.n85 4.5005
R8365 VOUT.n95 VOUT.n94 4.5005
R8366 VOUT.n104 VOUT.n103 4.5005
R8367 VOUT.n113 VOUT.n112 4.5005
R8368 VOUT.n122 VOUT.n121 4.5005
R8369 VOUT.n131 VOUT.n130 4.5005
R8370 VOUT.n140 VOUT.n139 4.5005
R8371 VOUT.n149 VOUT.n148 4.5005
R8372 VOUT.n158 VOUT.n157 4.5005
R8373 VOUT.n167 VOUT.n166 4.5005
R8374 VOUT.n176 VOUT.n175 4.5005
R8375 VOUT.n185 VOUT.n184 4.5005
R8376 VOUT.n1503 VOUT.n1502 4.14168
R8377 VOUT.n1494 VOUT.n1493 4.14168
R8378 VOUT.n1485 VOUT.n1484 4.14168
R8379 VOUT.n1476 VOUT.n1475 4.14168
R8380 VOUT.n1467 VOUT.n1466 4.14168
R8381 VOUT.n1458 VOUT.n1457 4.14168
R8382 VOUT.n1449 VOUT.n1448 4.14168
R8383 VOUT.n1440 VOUT.n1439 4.14168
R8384 VOUT.n1431 VOUT.n1430 4.14168
R8385 VOUT.n1422 VOUT.n1421 4.14168
R8386 VOUT.n1413 VOUT.n1412 4.14168
R8387 VOUT.n1404 VOUT.n1403 4.14168
R8388 VOUT.n1395 VOUT.n1394 4.14168
R8389 VOUT.n1386 VOUT.n1385 4.14168
R8390 VOUT.n1377 VOUT.n1376 4.14168
R8391 VOUT.n1368 VOUT.n1367 4.14168
R8392 VOUT.n1359 VOUT.n1358 4.14168
R8393 VOUT.n1350 VOUT.n1349 4.14168
R8394 VOUT.n1341 VOUT.n1340 4.14168
R8395 VOUT.n1332 VOUT.n1331 4.14168
R8396 VOUT.n1323 VOUT.n1322 4.14168
R8397 VOUT.n1127 VOUT.n1126 3.76521
R8398 VOUT.n1118 VOUT.n1117 3.76521
R8399 VOUT.n1109 VOUT.n1108 3.76521
R8400 VOUT.n1100 VOUT.n1099 3.76521
R8401 VOUT.n1091 VOUT.n1090 3.76521
R8402 VOUT.n1082 VOUT.n1081 3.76521
R8403 VOUT.n1073 VOUT.n1072 3.76521
R8404 VOUT.n1064 VOUT.n1063 3.76521
R8405 VOUT.n1055 VOUT.n1054 3.76521
R8406 VOUT.n1046 VOUT.n1045 3.76521
R8407 VOUT.n1037 VOUT.n1036 3.76521
R8408 VOUT.n1028 VOUT.n1027 3.76521
R8409 VOUT.n1019 VOUT.n1018 3.76521
R8410 VOUT.n1010 VOUT.n1009 3.76521
R8411 VOUT.n1001 VOUT.n1000 3.76521
R8412 VOUT.n992 VOUT.n991 3.76521
R8413 VOUT.n983 VOUT.n982 3.76521
R8414 VOUT.n974 VOUT.n973 3.76521
R8415 VOUT.n965 VOUT.n964 3.76521
R8416 VOUT.n956 VOUT.n955 3.76521
R8417 VOUT.n947 VOUT.n946 3.76521
R8418 VOUT.n1315 VOUT.n1314 3.76521
R8419 VOUT.n1306 VOUT.n1305 3.76521
R8420 VOUT.n1297 VOUT.n1296 3.76521
R8421 VOUT.n1288 VOUT.n1287 3.76521
R8422 VOUT.n1279 VOUT.n1278 3.76521
R8423 VOUT.n1270 VOUT.n1269 3.76521
R8424 VOUT.n1261 VOUT.n1260 3.76521
R8425 VOUT.n1252 VOUT.n1251 3.76521
R8426 VOUT.n1243 VOUT.n1242 3.76521
R8427 VOUT.n1234 VOUT.n1233 3.76521
R8428 VOUT.n1225 VOUT.n1224 3.76521
R8429 VOUT.n1216 VOUT.n1215 3.76521
R8430 VOUT.n1207 VOUT.n1206 3.76521
R8431 VOUT.n1198 VOUT.n1197 3.76521
R8432 VOUT.n1189 VOUT.n1188 3.76521
R8433 VOUT.n1180 VOUT.n1179 3.76521
R8434 VOUT.n1171 VOUT.n1170 3.76521
R8435 VOUT.n1162 VOUT.n1161 3.76521
R8436 VOUT.n1153 VOUT.n1152 3.76521
R8437 VOUT.n1144 VOUT.n1143 3.76521
R8438 VOUT.n1135 VOUT.n1134 3.76521
R8439 VOUT.n751 VOUT.n750 3.38874
R8440 VOUT.n742 VOUT.n741 3.38874
R8441 VOUT.n733 VOUT.n732 3.38874
R8442 VOUT.n724 VOUT.n723 3.38874
R8443 VOUT.n715 VOUT.n714 3.38874
R8444 VOUT.n706 VOUT.n705 3.38874
R8445 VOUT.n697 VOUT.n696 3.38874
R8446 VOUT.n688 VOUT.n687 3.38874
R8447 VOUT.n679 VOUT.n678 3.38874
R8448 VOUT.n670 VOUT.n669 3.38874
R8449 VOUT.n661 VOUT.n660 3.38874
R8450 VOUT.n652 VOUT.n651 3.38874
R8451 VOUT.n643 VOUT.n642 3.38874
R8452 VOUT.n634 VOUT.n633 3.38874
R8453 VOUT.n625 VOUT.n624 3.38874
R8454 VOUT.n616 VOUT.n615 3.38874
R8455 VOUT.n607 VOUT.n606 3.38874
R8456 VOUT.n598 VOUT.n597 3.38874
R8457 VOUT.n589 VOUT.n588 3.38874
R8458 VOUT.n580 VOUT.n579 3.38874
R8459 VOUT.n571 VOUT.n570 3.38874
R8460 VOUT.n939 VOUT.n938 3.38874
R8461 VOUT.n930 VOUT.n929 3.38874
R8462 VOUT.n921 VOUT.n920 3.38874
R8463 VOUT.n912 VOUT.n911 3.38874
R8464 VOUT.n903 VOUT.n902 3.38874
R8465 VOUT.n894 VOUT.n893 3.38874
R8466 VOUT.n885 VOUT.n884 3.38874
R8467 VOUT.n876 VOUT.n875 3.38874
R8468 VOUT.n867 VOUT.n866 3.38874
R8469 VOUT.n858 VOUT.n857 3.38874
R8470 VOUT.n849 VOUT.n848 3.38874
R8471 VOUT.n840 VOUT.n839 3.38874
R8472 VOUT.n831 VOUT.n830 3.38874
R8473 VOUT.n822 VOUT.n821 3.38874
R8474 VOUT.n813 VOUT.n812 3.38874
R8475 VOUT.n804 VOUT.n803 3.38874
R8476 VOUT.n795 VOUT.n794 3.38874
R8477 VOUT.n786 VOUT.n785 3.38874
R8478 VOUT.n777 VOUT.n776 3.38874
R8479 VOUT.n768 VOUT.n767 3.38874
R8480 VOUT.n759 VOUT.n758 3.38874
R8481 VOUT.n2067 VOUT.n2066 3.38874
R8482 VOUT.n2058 VOUT.n2057 3.38874
R8483 VOUT.n2049 VOUT.n2048 3.38874
R8484 VOUT.n2040 VOUT.n2039 3.38874
R8485 VOUT.n2031 VOUT.n2030 3.38874
R8486 VOUT.n2022 VOUT.n2021 3.38874
R8487 VOUT.n2013 VOUT.n2012 3.38874
R8488 VOUT.n2004 VOUT.n2003 3.38874
R8489 VOUT.n1995 VOUT.n1994 3.38874
R8490 VOUT.n1986 VOUT.n1985 3.38874
R8491 VOUT.n1977 VOUT.n1976 3.38874
R8492 VOUT.n1968 VOUT.n1967 3.38874
R8493 VOUT.n1959 VOUT.n1958 3.38874
R8494 VOUT.n1950 VOUT.n1949 3.38874
R8495 VOUT.n1941 VOUT.n1940 3.38874
R8496 VOUT.n1932 VOUT.n1931 3.38874
R8497 VOUT.n1923 VOUT.n1922 3.38874
R8498 VOUT.n1914 VOUT.n1913 3.38874
R8499 VOUT.n1905 VOUT.n1904 3.38874
R8500 VOUT.n1896 VOUT.n1895 3.38874
R8501 VOUT.n1887 VOUT.n1886 3.38874
R8502 VOUT.n572 VOUT.n571 3.02889
R8503 VOUT.n581 VOUT.n580 3.02889
R8504 VOUT.n590 VOUT.n589 3.02889
R8505 VOUT.n599 VOUT.n598 3.02889
R8506 VOUT.n608 VOUT.n607 3.02889
R8507 VOUT.n617 VOUT.n616 3.02889
R8508 VOUT.n626 VOUT.n625 3.02889
R8509 VOUT.n635 VOUT.n634 3.02889
R8510 VOUT.n644 VOUT.n643 3.02889
R8511 VOUT.n653 VOUT.n652 3.02889
R8512 VOUT.n662 VOUT.n661 3.02889
R8513 VOUT.n671 VOUT.n670 3.02889
R8514 VOUT.n680 VOUT.n679 3.02889
R8515 VOUT.n689 VOUT.n688 3.02889
R8516 VOUT.n698 VOUT.n697 3.02889
R8517 VOUT.n707 VOUT.n706 3.02889
R8518 VOUT.n716 VOUT.n715 3.02889
R8519 VOUT.n725 VOUT.n724 3.02889
R8520 VOUT.n734 VOUT.n733 3.02889
R8521 VOUT.n743 VOUT.n742 3.02889
R8522 VOUT.n752 VOUT.n751 3.02889
R8523 VOUT.n760 VOUT.n759 3.02889
R8524 VOUT.n769 VOUT.n768 3.02889
R8525 VOUT.n778 VOUT.n777 3.02889
R8526 VOUT.n787 VOUT.n786 3.02889
R8527 VOUT.n796 VOUT.n795 3.02889
R8528 VOUT.n805 VOUT.n804 3.02889
R8529 VOUT.n814 VOUT.n813 3.02889
R8530 VOUT.n823 VOUT.n822 3.02889
R8531 VOUT.n832 VOUT.n831 3.02889
R8532 VOUT.n841 VOUT.n840 3.02889
R8533 VOUT.n850 VOUT.n849 3.02889
R8534 VOUT.n859 VOUT.n858 3.02889
R8535 VOUT.n868 VOUT.n867 3.02889
R8536 VOUT.n877 VOUT.n876 3.02889
R8537 VOUT.n886 VOUT.n885 3.02889
R8538 VOUT.n895 VOUT.n894 3.02889
R8539 VOUT.n904 VOUT.n903 3.02889
R8540 VOUT.n913 VOUT.n912 3.02889
R8541 VOUT.n922 VOUT.n921 3.02889
R8542 VOUT.n931 VOUT.n930 3.02889
R8543 VOUT.n940 VOUT.n939 3.02889
R8544 VOUT.n948 VOUT.n947 3.02889
R8545 VOUT.n957 VOUT.n956 3.02889
R8546 VOUT.n966 VOUT.n965 3.02889
R8547 VOUT.n975 VOUT.n974 3.02889
R8548 VOUT.n984 VOUT.n983 3.02889
R8549 VOUT.n993 VOUT.n992 3.02889
R8550 VOUT.n1002 VOUT.n1001 3.02889
R8551 VOUT.n1011 VOUT.n1010 3.02889
R8552 VOUT.n1020 VOUT.n1019 3.02889
R8553 VOUT.n1029 VOUT.n1028 3.02889
R8554 VOUT.n1038 VOUT.n1037 3.02889
R8555 VOUT.n1047 VOUT.n1046 3.02889
R8556 VOUT.n1056 VOUT.n1055 3.02889
R8557 VOUT.n1065 VOUT.n1064 3.02889
R8558 VOUT.n1074 VOUT.n1073 3.02889
R8559 VOUT.n1083 VOUT.n1082 3.02889
R8560 VOUT.n1092 VOUT.n1091 3.02889
R8561 VOUT.n1101 VOUT.n1100 3.02889
R8562 VOUT.n1110 VOUT.n1109 3.02889
R8563 VOUT.n1119 VOUT.n1118 3.02889
R8564 VOUT.n1128 VOUT.n1127 3.02889
R8565 VOUT.n1136 VOUT.n1135 3.02889
R8566 VOUT.n1145 VOUT.n1144 3.02889
R8567 VOUT.n1154 VOUT.n1153 3.02889
R8568 VOUT.n1163 VOUT.n1162 3.02889
R8569 VOUT.n1172 VOUT.n1171 3.02889
R8570 VOUT.n1181 VOUT.n1180 3.02889
R8571 VOUT.n1190 VOUT.n1189 3.02889
R8572 VOUT.n1199 VOUT.n1198 3.02889
R8573 VOUT.n1208 VOUT.n1207 3.02889
R8574 VOUT.n1217 VOUT.n1216 3.02889
R8575 VOUT.n1226 VOUT.n1225 3.02889
R8576 VOUT.n1235 VOUT.n1234 3.02889
R8577 VOUT.n1244 VOUT.n1243 3.02889
R8578 VOUT.n1253 VOUT.n1252 3.02889
R8579 VOUT.n1262 VOUT.n1261 3.02889
R8580 VOUT.n1271 VOUT.n1270 3.02889
R8581 VOUT.n1280 VOUT.n1279 3.02889
R8582 VOUT.n1289 VOUT.n1288 3.02889
R8583 VOUT.n1298 VOUT.n1297 3.02889
R8584 VOUT.n1307 VOUT.n1306 3.02889
R8585 VOUT.n1316 VOUT.n1315 3.02889
R8586 VOUT.n1324 VOUT.n1323 3.02889
R8587 VOUT.n1333 VOUT.n1332 3.02889
R8588 VOUT.n1342 VOUT.n1341 3.02889
R8589 VOUT.n1351 VOUT.n1350 3.02889
R8590 VOUT.n1360 VOUT.n1359 3.02889
R8591 VOUT.n1369 VOUT.n1368 3.02889
R8592 VOUT.n1378 VOUT.n1377 3.02889
R8593 VOUT.n1387 VOUT.n1386 3.02889
R8594 VOUT.n1396 VOUT.n1395 3.02889
R8595 VOUT.n1405 VOUT.n1404 3.02889
R8596 VOUT.n1414 VOUT.n1413 3.02889
R8597 VOUT.n1423 VOUT.n1422 3.02889
R8598 VOUT.n1432 VOUT.n1431 3.02889
R8599 VOUT.n1441 VOUT.n1440 3.02889
R8600 VOUT.n1450 VOUT.n1449 3.02889
R8601 VOUT.n1459 VOUT.n1458 3.02889
R8602 VOUT.n1468 VOUT.n1467 3.02889
R8603 VOUT.n1477 VOUT.n1476 3.02889
R8604 VOUT.n1486 VOUT.n1485 3.02889
R8605 VOUT.n1495 VOUT.n1494 3.02889
R8606 VOUT.n1504 VOUT.n1503 3.02889
R8607 VOUT.n1512 VOUT.n1511 3.02889
R8608 VOUT.n1521 VOUT.n1520 3.02889
R8609 VOUT.n1530 VOUT.n1529 3.02889
R8610 VOUT.n1539 VOUT.n1538 3.02889
R8611 VOUT.n1548 VOUT.n1547 3.02889
R8612 VOUT.n1557 VOUT.n1556 3.02889
R8613 VOUT.n1566 VOUT.n1565 3.02889
R8614 VOUT.n1575 VOUT.n1574 3.02889
R8615 VOUT.n1584 VOUT.n1583 3.02889
R8616 VOUT.n1593 VOUT.n1592 3.02889
R8617 VOUT.n1602 VOUT.n1601 3.02889
R8618 VOUT.n1611 VOUT.n1610 3.02889
R8619 VOUT.n1620 VOUT.n1619 3.02889
R8620 VOUT.n1629 VOUT.n1628 3.02889
R8621 VOUT.n1638 VOUT.n1637 3.02889
R8622 VOUT.n1647 VOUT.n1646 3.02889
R8623 VOUT.n1656 VOUT.n1655 3.02889
R8624 VOUT.n1665 VOUT.n1664 3.02889
R8625 VOUT.n1674 VOUT.n1673 3.02889
R8626 VOUT.n1683 VOUT.n1682 3.02889
R8627 VOUT.n1692 VOUT.n1691 3.02889
R8628 VOUT.n1700 VOUT.n1699 3.02889
R8629 VOUT.n1709 VOUT.n1708 3.02889
R8630 VOUT.n1718 VOUT.n1717 3.02889
R8631 VOUT.n1727 VOUT.n1726 3.02889
R8632 VOUT.n1736 VOUT.n1735 3.02889
R8633 VOUT.n1745 VOUT.n1744 3.02889
R8634 VOUT.n1754 VOUT.n1753 3.02889
R8635 VOUT.n1763 VOUT.n1762 3.02889
R8636 VOUT.n1772 VOUT.n1771 3.02889
R8637 VOUT.n1781 VOUT.n1780 3.02889
R8638 VOUT.n1790 VOUT.n1789 3.02889
R8639 VOUT.n1799 VOUT.n1798 3.02889
R8640 VOUT.n1808 VOUT.n1807 3.02889
R8641 VOUT.n1817 VOUT.n1816 3.02889
R8642 VOUT.n1826 VOUT.n1825 3.02889
R8643 VOUT.n1835 VOUT.n1834 3.02889
R8644 VOUT.n1844 VOUT.n1843 3.02889
R8645 VOUT.n1853 VOUT.n1852 3.02889
R8646 VOUT.n1862 VOUT.n1861 3.02889
R8647 VOUT.n1871 VOUT.n1870 3.02889
R8648 VOUT.n1880 VOUT.n1879 3.02889
R8649 VOUT.n1888 VOUT.n1887 3.02889
R8650 VOUT.n1897 VOUT.n1896 3.02889
R8651 VOUT.n1906 VOUT.n1905 3.02889
R8652 VOUT.n1915 VOUT.n1914 3.02889
R8653 VOUT.n1924 VOUT.n1923 3.02889
R8654 VOUT.n1933 VOUT.n1932 3.02889
R8655 VOUT.n1942 VOUT.n1941 3.02889
R8656 VOUT.n1951 VOUT.n1950 3.02889
R8657 VOUT.n1960 VOUT.n1959 3.02889
R8658 VOUT.n1969 VOUT.n1968 3.02889
R8659 VOUT.n1978 VOUT.n1977 3.02889
R8660 VOUT.n1987 VOUT.n1986 3.02889
R8661 VOUT.n1996 VOUT.n1995 3.02889
R8662 VOUT.n2005 VOUT.n2004 3.02889
R8663 VOUT.n2014 VOUT.n2013 3.02889
R8664 VOUT.n2023 VOUT.n2022 3.02889
R8665 VOUT.n2032 VOUT.n2031 3.02889
R8666 VOUT.n2041 VOUT.n2040 3.02889
R8667 VOUT.n2050 VOUT.n2049 3.02889
R8668 VOUT.n2059 VOUT.n2058 3.02889
R8669 VOUT.n2068 VOUT.n2067 3.02889
R8670 VOUT.n2076 VOUT.n2075 3.02889
R8671 VOUT.n2085 VOUT.n2084 3.02889
R8672 VOUT.n2094 VOUT.n2093 3.02889
R8673 VOUT.n2103 VOUT.n2102 3.02889
R8674 VOUT.n2112 VOUT.n2111 3.02889
R8675 VOUT.n2121 VOUT.n2120 3.02889
R8676 VOUT.n2130 VOUT.n2129 3.02889
R8677 VOUT.n2139 VOUT.n2138 3.02889
R8678 VOUT.n2148 VOUT.n2147 3.02889
R8679 VOUT.n2157 VOUT.n2156 3.02889
R8680 VOUT.n2166 VOUT.n2165 3.02889
R8681 VOUT.n2175 VOUT.n2174 3.02889
R8682 VOUT.n2184 VOUT.n2183 3.02889
R8683 VOUT.n2193 VOUT.n2192 3.02889
R8684 VOUT.n2202 VOUT.n2201 3.02889
R8685 VOUT.n2211 VOUT.n2210 3.02889
R8686 VOUT.n2220 VOUT.n2219 3.02889
R8687 VOUT.n2229 VOUT.n2228 3.02889
R8688 VOUT.n2238 VOUT.n2237 3.02889
R8689 VOUT.n2247 VOUT.n2246 3.02889
R8690 VOUT.n2256 VOUT.n2255 3.02889
R8691 VOUT.n2397 VOUT.n2396 3.02889
R8692 VOUT.n2390 VOUT.n2389 3.02889
R8693 VOUT.n2383 VOUT.n2382 3.02889
R8694 VOUT.n2376 VOUT.n2375 3.02889
R8695 VOUT.n2369 VOUT.n2368 3.02889
R8696 VOUT.n2362 VOUT.n2361 3.02889
R8697 VOUT.n2355 VOUT.n2354 3.02889
R8698 VOUT.n2348 VOUT.n2347 3.02889
R8699 VOUT.n2341 VOUT.n2340 3.02889
R8700 VOUT.n2334 VOUT.n2333 3.02889
R8701 VOUT.n2327 VOUT.n2326 3.02889
R8702 VOUT.n2320 VOUT.n2319 3.02889
R8703 VOUT.n2313 VOUT.n2312 3.02889
R8704 VOUT.n2306 VOUT.n2305 3.02889
R8705 VOUT.n2299 VOUT.n2298 3.02889
R8706 VOUT.n2292 VOUT.n2291 3.02889
R8707 VOUT.n2285 VOUT.n2284 3.02889
R8708 VOUT.n2278 VOUT.n2277 3.02889
R8709 VOUT.n2271 VOUT.n2270 3.02889
R8710 VOUT.n2264 VOUT.n2263 3.02889
R8711 VOUT.n2404 VOUT.n2403 3.02889
R8712 VOUT.n1879 VOUT.n1878 3.01226
R8713 VOUT.n1870 VOUT.n1869 3.01226
R8714 VOUT.n1861 VOUT.n1860 3.01226
R8715 VOUT.n1852 VOUT.n1851 3.01226
R8716 VOUT.n1843 VOUT.n1842 3.01226
R8717 VOUT.n1834 VOUT.n1833 3.01226
R8718 VOUT.n1825 VOUT.n1824 3.01226
R8719 VOUT.n1816 VOUT.n1815 3.01226
R8720 VOUT.n1807 VOUT.n1806 3.01226
R8721 VOUT.n1798 VOUT.n1797 3.01226
R8722 VOUT.n1789 VOUT.n1788 3.01226
R8723 VOUT.n1780 VOUT.n1779 3.01226
R8724 VOUT.n1771 VOUT.n1770 3.01226
R8725 VOUT.n1762 VOUT.n1761 3.01226
R8726 VOUT.n1753 VOUT.n1752 3.01226
R8727 VOUT.n1744 VOUT.n1743 3.01226
R8728 VOUT.n1735 VOUT.n1734 3.01226
R8729 VOUT.n1726 VOUT.n1725 3.01226
R8730 VOUT.n1717 VOUT.n1716 3.01226
R8731 VOUT.n1708 VOUT.n1707 3.01226
R8732 VOUT.n1699 VOUT.n1698 3.01226
R8733 VOUT.n2255 VOUT.n2254 2.63579
R8734 VOUT.n2246 VOUT.n2245 2.63579
R8735 VOUT.n2237 VOUT.n2236 2.63579
R8736 VOUT.n2228 VOUT.n2227 2.63579
R8737 VOUT.n2219 VOUT.n2218 2.63579
R8738 VOUT.n2210 VOUT.n2209 2.63579
R8739 VOUT.n2201 VOUT.n2200 2.63579
R8740 VOUT.n2192 VOUT.n2191 2.63579
R8741 VOUT.n2183 VOUT.n2182 2.63579
R8742 VOUT.n2174 VOUT.n2173 2.63579
R8743 VOUT.n2165 VOUT.n2164 2.63579
R8744 VOUT.n2156 VOUT.n2155 2.63579
R8745 VOUT.n2147 VOUT.n2146 2.63579
R8746 VOUT.n2138 VOUT.n2137 2.63579
R8747 VOUT.n2129 VOUT.n2128 2.63579
R8748 VOUT.n2120 VOUT.n2119 2.63579
R8749 VOUT.n2111 VOUT.n2110 2.63579
R8750 VOUT.n2102 VOUT.n2101 2.63579
R8751 VOUT.n2093 VOUT.n2092 2.63579
R8752 VOUT.n2084 VOUT.n2083 2.63579
R8753 VOUT.n2075 VOUT.n2074 2.63579
R8754 VOUT.n560 VOUT.n559 2.63579
R8755 VOUT.n551 VOUT.n550 2.63579
R8756 VOUT.n542 VOUT.n541 2.63579
R8757 VOUT.n533 VOUT.n532 2.63579
R8758 VOUT.n524 VOUT.n523 2.63579
R8759 VOUT.n515 VOUT.n514 2.63579
R8760 VOUT.n506 VOUT.n505 2.63579
R8761 VOUT.n497 VOUT.n496 2.63579
R8762 VOUT.n488 VOUT.n487 2.63579
R8763 VOUT.n479 VOUT.n478 2.63579
R8764 VOUT.n470 VOUT.n469 2.63579
R8765 VOUT.n461 VOUT.n460 2.63579
R8766 VOUT.n452 VOUT.n451 2.63579
R8767 VOUT.n443 VOUT.n442 2.63579
R8768 VOUT.n434 VOUT.n433 2.63579
R8769 VOUT.n425 VOUT.n424 2.63579
R8770 VOUT.n416 VOUT.n415 2.63579
R8771 VOUT.n407 VOUT.n406 2.63579
R8772 VOUT.n398 VOUT.n397 2.63579
R8773 VOUT.n389 VOUT.n388 2.63579
R8774 VOUT.n381 VOUT.n380 2.63579
R8775 VOUT.n372 VOUT.n371 2.63579
R8776 VOUT.n363 VOUT.n362 2.63579
R8777 VOUT.n354 VOUT.n353 2.63579
R8778 VOUT.n345 VOUT.n344 2.63579
R8779 VOUT.n336 VOUT.n335 2.63579
R8780 VOUT.n327 VOUT.n326 2.63579
R8781 VOUT.n318 VOUT.n317 2.63579
R8782 VOUT.n309 VOUT.n308 2.63579
R8783 VOUT.n300 VOUT.n299 2.63579
R8784 VOUT.n291 VOUT.n290 2.63579
R8785 VOUT.n282 VOUT.n281 2.63579
R8786 VOUT.n273 VOUT.n272 2.63579
R8787 VOUT.n264 VOUT.n263 2.63579
R8788 VOUT.n255 VOUT.n254 2.63579
R8789 VOUT.n246 VOUT.n245 2.63579
R8790 VOUT.n237 VOUT.n236 2.63579
R8791 VOUT.n228 VOUT.n227 2.63579
R8792 VOUT.n219 VOUT.n218 2.63579
R8793 VOUT.n210 VOUT.n209 2.63579
R8794 VOUT.n201 VOUT.n200 2.63579
R8795 VOUT.n193 VOUT.n192 2.63579
R8796 VOUT.n184 VOUT.n183 2.63579
R8797 VOUT.n175 VOUT.n174 2.63579
R8798 VOUT.n166 VOUT.n165 2.63579
R8799 VOUT.n157 VOUT.n156 2.63579
R8800 VOUT.n148 VOUT.n147 2.63579
R8801 VOUT.n139 VOUT.n138 2.63579
R8802 VOUT.n130 VOUT.n129 2.63579
R8803 VOUT.n121 VOUT.n120 2.63579
R8804 VOUT.n112 VOUT.n111 2.63579
R8805 VOUT.n103 VOUT.n102 2.63579
R8806 VOUT.n94 VOUT.n93 2.63579
R8807 VOUT.n85 VOUT.n84 2.63579
R8808 VOUT.n76 VOUT.n75 2.63579
R8809 VOUT.n67 VOUT.n66 2.63579
R8810 VOUT.n58 VOUT.n57 2.63579
R8811 VOUT.n49 VOUT.n48 2.63579
R8812 VOUT.n40 VOUT.n39 2.63579
R8813 VOUT.n31 VOUT.n30 2.63579
R8814 VOUT.n22 VOUT.n21 2.63579
R8815 VOUT.n13 VOUT.n12 2.63579
R8816 VOUT.n5 VOUT.n4 2.63579
R8817 VOUT.n2263 VOUT.n2262 1.88285
R8818 VOUT.n2270 VOUT.n2269 1.88285
R8819 VOUT.n2277 VOUT.n2276 1.88285
R8820 VOUT.n2284 VOUT.n2283 1.88285
R8821 VOUT.n2291 VOUT.n2290 1.88285
R8822 VOUT.n2298 VOUT.n2297 1.88285
R8823 VOUT.n2305 VOUT.n2304 1.88285
R8824 VOUT.n2312 VOUT.n2311 1.88285
R8825 VOUT.n2319 VOUT.n2318 1.88285
R8826 VOUT.n2326 VOUT.n2325 1.88285
R8827 VOUT.n2333 VOUT.n2332 1.88285
R8828 VOUT.n2340 VOUT.n2339 1.88285
R8829 VOUT.n2347 VOUT.n2346 1.88285
R8830 VOUT.n2354 VOUT.n2353 1.88285
R8831 VOUT.n2361 VOUT.n2360 1.88285
R8832 VOUT.n2368 VOUT.n2367 1.88285
R8833 VOUT.n2375 VOUT.n2374 1.88285
R8834 VOUT.n2382 VOUT.n2381 1.88285
R8835 VOUT.n2389 VOUT.n2388 1.88285
R8836 VOUT.n2396 VOUT.n2395 1.88285
R8837 VOUT.n2403 VOUT.n2402 1.88285
R8838 VOUT.n383 VOUT.n382 1.19441
R8839 VOUT.n195 VOUT.n194 1.19441
R8840 VOUT.n7 VOUT.n6 1.19441
R8841 VOUT.n2445 VOUT.n2264 1.15278
R8842 VOUT.n2443 VOUT.n2271 1.15278
R8843 VOUT.n2441 VOUT.n2278 1.15278
R8844 VOUT.n2439 VOUT.n2285 1.15278
R8845 VOUT.n2437 VOUT.n2292 1.15278
R8846 VOUT.n2435 VOUT.n2299 1.15278
R8847 VOUT.n2433 VOUT.n2306 1.15278
R8848 VOUT.n2431 VOUT.n2313 1.15278
R8849 VOUT.n2429 VOUT.n2320 1.15278
R8850 VOUT.n2427 VOUT.n2327 1.15278
R8851 VOUT.n2425 VOUT.n2334 1.15278
R8852 VOUT.n2423 VOUT.n2341 1.15278
R8853 VOUT.n2421 VOUT.n2348 1.15278
R8854 VOUT.n2419 VOUT.n2355 1.15278
R8855 VOUT.n2417 VOUT.n2362 1.15278
R8856 VOUT.n2415 VOUT.n2369 1.15278
R8857 VOUT.n2413 VOUT.n2376 1.15278
R8858 VOUT.n2411 VOUT.n2383 1.15278
R8859 VOUT.n2409 VOUT.n2390 1.15278
R8860 VOUT.n2407 VOUT.n2397 1.15278
R8861 VOUT.n753 VOUT.n752 1.15278
R8862 VOUT.n744 VOUT.n743 1.15278
R8863 VOUT.n735 VOUT.n734 1.15278
R8864 VOUT.n726 VOUT.n725 1.15278
R8865 VOUT.n717 VOUT.n716 1.15278
R8866 VOUT.n708 VOUT.n707 1.15278
R8867 VOUT.n699 VOUT.n698 1.15278
R8868 VOUT.n690 VOUT.n689 1.15278
R8869 VOUT.n681 VOUT.n680 1.15278
R8870 VOUT.n672 VOUT.n671 1.15278
R8871 VOUT.n663 VOUT.n662 1.15278
R8872 VOUT.n654 VOUT.n653 1.15278
R8873 VOUT.n645 VOUT.n644 1.15278
R8874 VOUT.n636 VOUT.n635 1.15278
R8875 VOUT.n627 VOUT.n626 1.15278
R8876 VOUT.n618 VOUT.n617 1.15278
R8877 VOUT.n609 VOUT.n608 1.15278
R8878 VOUT.n600 VOUT.n599 1.15278
R8879 VOUT.n591 VOUT.n590 1.15278
R8880 VOUT.n582 VOUT.n581 1.15278
R8881 VOUT.n573 VOUT.n572 1.15278
R8882 VOUT.n941 VOUT.n940 1.15278
R8883 VOUT.n932 VOUT.n931 1.15278
R8884 VOUT.n923 VOUT.n922 1.15278
R8885 VOUT.n914 VOUT.n913 1.15278
R8886 VOUT.n905 VOUT.n904 1.15278
R8887 VOUT.n896 VOUT.n895 1.15278
R8888 VOUT.n887 VOUT.n886 1.15278
R8889 VOUT.n878 VOUT.n877 1.15278
R8890 VOUT.n869 VOUT.n868 1.15278
R8891 VOUT.n860 VOUT.n859 1.15278
R8892 VOUT.n851 VOUT.n850 1.15278
R8893 VOUT.n842 VOUT.n841 1.15278
R8894 VOUT.n833 VOUT.n832 1.15278
R8895 VOUT.n824 VOUT.n823 1.15278
R8896 VOUT.n815 VOUT.n814 1.15278
R8897 VOUT.n806 VOUT.n805 1.15278
R8898 VOUT.n797 VOUT.n796 1.15278
R8899 VOUT.n788 VOUT.n787 1.15278
R8900 VOUT.n779 VOUT.n778 1.15278
R8901 VOUT.n770 VOUT.n769 1.15278
R8902 VOUT.n761 VOUT.n760 1.15278
R8903 VOUT.n1129 VOUT.n1128 1.15278
R8904 VOUT.n1120 VOUT.n1119 1.15278
R8905 VOUT.n1111 VOUT.n1110 1.15278
R8906 VOUT.n1102 VOUT.n1101 1.15278
R8907 VOUT.n1093 VOUT.n1092 1.15278
R8908 VOUT.n1084 VOUT.n1083 1.15278
R8909 VOUT.n1075 VOUT.n1074 1.15278
R8910 VOUT.n1066 VOUT.n1065 1.15278
R8911 VOUT.n1057 VOUT.n1056 1.15278
R8912 VOUT.n1048 VOUT.n1047 1.15278
R8913 VOUT.n1039 VOUT.n1038 1.15278
R8914 VOUT.n1030 VOUT.n1029 1.15278
R8915 VOUT.n1021 VOUT.n1020 1.15278
R8916 VOUT.n1012 VOUT.n1011 1.15278
R8917 VOUT.n1003 VOUT.n1002 1.15278
R8918 VOUT.n994 VOUT.n993 1.15278
R8919 VOUT.n985 VOUT.n984 1.15278
R8920 VOUT.n976 VOUT.n975 1.15278
R8921 VOUT.n967 VOUT.n966 1.15278
R8922 VOUT.n958 VOUT.n957 1.15278
R8923 VOUT.n949 VOUT.n948 1.15278
R8924 VOUT.n1317 VOUT.n1316 1.15278
R8925 VOUT.n1308 VOUT.n1307 1.15278
R8926 VOUT.n1299 VOUT.n1298 1.15278
R8927 VOUT.n1290 VOUT.n1289 1.15278
R8928 VOUT.n1281 VOUT.n1280 1.15278
R8929 VOUT.n1272 VOUT.n1271 1.15278
R8930 VOUT.n1263 VOUT.n1262 1.15278
R8931 VOUT.n1254 VOUT.n1253 1.15278
R8932 VOUT.n1245 VOUT.n1244 1.15278
R8933 VOUT.n1236 VOUT.n1235 1.15278
R8934 VOUT.n1227 VOUT.n1226 1.15278
R8935 VOUT.n1218 VOUT.n1217 1.15278
R8936 VOUT.n1209 VOUT.n1208 1.15278
R8937 VOUT.n1200 VOUT.n1199 1.15278
R8938 VOUT.n1191 VOUT.n1190 1.15278
R8939 VOUT.n1182 VOUT.n1181 1.15278
R8940 VOUT.n1173 VOUT.n1172 1.15278
R8941 VOUT.n1164 VOUT.n1163 1.15278
R8942 VOUT.n1155 VOUT.n1154 1.15278
R8943 VOUT.n1146 VOUT.n1145 1.15278
R8944 VOUT.n1137 VOUT.n1136 1.15278
R8945 VOUT.n1505 VOUT.n1504 1.15278
R8946 VOUT.n1496 VOUT.n1495 1.15278
R8947 VOUT.n1487 VOUT.n1486 1.15278
R8948 VOUT.n1478 VOUT.n1477 1.15278
R8949 VOUT.n1469 VOUT.n1468 1.15278
R8950 VOUT.n1460 VOUT.n1459 1.15278
R8951 VOUT.n1451 VOUT.n1450 1.15278
R8952 VOUT.n1442 VOUT.n1441 1.15278
R8953 VOUT.n1433 VOUT.n1432 1.15278
R8954 VOUT.n1424 VOUT.n1423 1.15278
R8955 VOUT.n1415 VOUT.n1414 1.15278
R8956 VOUT.n1406 VOUT.n1405 1.15278
R8957 VOUT.n1397 VOUT.n1396 1.15278
R8958 VOUT.n1388 VOUT.n1387 1.15278
R8959 VOUT.n1379 VOUT.n1378 1.15278
R8960 VOUT.n1370 VOUT.n1369 1.15278
R8961 VOUT.n1361 VOUT.n1360 1.15278
R8962 VOUT.n1352 VOUT.n1351 1.15278
R8963 VOUT.n1343 VOUT.n1342 1.15278
R8964 VOUT.n1334 VOUT.n1333 1.15278
R8965 VOUT.n1325 VOUT.n1324 1.15278
R8966 VOUT.n1693 VOUT.n1692 1.15278
R8967 VOUT.n1684 VOUT.n1683 1.15278
R8968 VOUT.n1675 VOUT.n1674 1.15278
R8969 VOUT.n1666 VOUT.n1665 1.15278
R8970 VOUT.n1657 VOUT.n1656 1.15278
R8971 VOUT.n1648 VOUT.n1647 1.15278
R8972 VOUT.n1639 VOUT.n1638 1.15278
R8973 VOUT.n1630 VOUT.n1629 1.15278
R8974 VOUT.n1621 VOUT.n1620 1.15278
R8975 VOUT.n1612 VOUT.n1611 1.15278
R8976 VOUT.n1603 VOUT.n1602 1.15278
R8977 VOUT.n1594 VOUT.n1593 1.15278
R8978 VOUT.n1585 VOUT.n1584 1.15278
R8979 VOUT.n1576 VOUT.n1575 1.15278
R8980 VOUT.n1567 VOUT.n1566 1.15278
R8981 VOUT.n1558 VOUT.n1557 1.15278
R8982 VOUT.n1549 VOUT.n1548 1.15278
R8983 VOUT.n1540 VOUT.n1539 1.15278
R8984 VOUT.n1531 VOUT.n1530 1.15278
R8985 VOUT.n1522 VOUT.n1521 1.15278
R8986 VOUT.n1513 VOUT.n1512 1.15278
R8987 VOUT.n1881 VOUT.n1880 1.15278
R8988 VOUT.n1872 VOUT.n1871 1.15278
R8989 VOUT.n1863 VOUT.n1862 1.15278
R8990 VOUT.n1854 VOUT.n1853 1.15278
R8991 VOUT.n1845 VOUT.n1844 1.15278
R8992 VOUT.n1836 VOUT.n1835 1.15278
R8993 VOUT.n1827 VOUT.n1826 1.15278
R8994 VOUT.n1818 VOUT.n1817 1.15278
R8995 VOUT.n1809 VOUT.n1808 1.15278
R8996 VOUT.n1800 VOUT.n1799 1.15278
R8997 VOUT.n1791 VOUT.n1790 1.15278
R8998 VOUT.n1782 VOUT.n1781 1.15278
R8999 VOUT.n1773 VOUT.n1772 1.15278
R9000 VOUT.n1764 VOUT.n1763 1.15278
R9001 VOUT.n1755 VOUT.n1754 1.15278
R9002 VOUT.n1746 VOUT.n1745 1.15278
R9003 VOUT.n1737 VOUT.n1736 1.15278
R9004 VOUT.n1728 VOUT.n1727 1.15278
R9005 VOUT.n1719 VOUT.n1718 1.15278
R9006 VOUT.n1710 VOUT.n1709 1.15278
R9007 VOUT.n1701 VOUT.n1700 1.15278
R9008 VOUT.n2069 VOUT.n2068 1.15278
R9009 VOUT.n2060 VOUT.n2059 1.15278
R9010 VOUT.n2051 VOUT.n2050 1.15278
R9011 VOUT.n2042 VOUT.n2041 1.15278
R9012 VOUT.n2033 VOUT.n2032 1.15278
R9013 VOUT.n2024 VOUT.n2023 1.15278
R9014 VOUT.n2015 VOUT.n2014 1.15278
R9015 VOUT.n2006 VOUT.n2005 1.15278
R9016 VOUT.n1997 VOUT.n1996 1.15278
R9017 VOUT.n1988 VOUT.n1987 1.15278
R9018 VOUT.n1979 VOUT.n1978 1.15278
R9019 VOUT.n1970 VOUT.n1969 1.15278
R9020 VOUT.n1961 VOUT.n1960 1.15278
R9021 VOUT.n1952 VOUT.n1951 1.15278
R9022 VOUT.n1943 VOUT.n1942 1.15278
R9023 VOUT.n1934 VOUT.n1933 1.15278
R9024 VOUT.n1925 VOUT.n1924 1.15278
R9025 VOUT.n1916 VOUT.n1915 1.15278
R9026 VOUT.n1907 VOUT.n1906 1.15278
R9027 VOUT.n1898 VOUT.n1897 1.15278
R9028 VOUT.n1889 VOUT.n1888 1.15278
R9029 VOUT.n2257 VOUT.n2256 1.15278
R9030 VOUT.n2248 VOUT.n2247 1.15278
R9031 VOUT.n2239 VOUT.n2238 1.15278
R9032 VOUT.n2230 VOUT.n2229 1.15278
R9033 VOUT.n2221 VOUT.n2220 1.15278
R9034 VOUT.n2212 VOUT.n2211 1.15278
R9035 VOUT.n2203 VOUT.n2202 1.15278
R9036 VOUT.n2194 VOUT.n2193 1.15278
R9037 VOUT.n2185 VOUT.n2184 1.15278
R9038 VOUT.n2176 VOUT.n2175 1.15278
R9039 VOUT.n2167 VOUT.n2166 1.15278
R9040 VOUT.n2158 VOUT.n2157 1.15278
R9041 VOUT.n2149 VOUT.n2148 1.15278
R9042 VOUT.n2140 VOUT.n2139 1.15278
R9043 VOUT.n2131 VOUT.n2130 1.15278
R9044 VOUT.n2122 VOUT.n2121 1.15278
R9045 VOUT.n2113 VOUT.n2112 1.15278
R9046 VOUT.n2104 VOUT.n2103 1.15278
R9047 VOUT.n2095 VOUT.n2094 1.15278
R9048 VOUT.n2086 VOUT.n2085 1.15278
R9049 VOUT.n2077 VOUT.n2076 1.15278
R9050 VOUT.n2405 VOUT.n2404 1.15278
R9051 VOUT.n391 VOUT.n390 1.13663
R9052 VOUT.n400 VOUT.n399 1.13663
R9053 VOUT.n409 VOUT.n408 1.13663
R9054 VOUT.n418 VOUT.n417 1.13663
R9055 VOUT.n427 VOUT.n426 1.13663
R9056 VOUT.n436 VOUT.n435 1.13663
R9057 VOUT.n445 VOUT.n444 1.13663
R9058 VOUT.n454 VOUT.n453 1.13663
R9059 VOUT.n463 VOUT.n462 1.13663
R9060 VOUT.n472 VOUT.n471 1.13663
R9061 VOUT.n481 VOUT.n480 1.13663
R9062 VOUT.n490 VOUT.n489 1.13663
R9063 VOUT.n499 VOUT.n498 1.13663
R9064 VOUT.n508 VOUT.n507 1.13663
R9065 VOUT.n517 VOUT.n516 1.13663
R9066 VOUT.n526 VOUT.n525 1.13663
R9067 VOUT.n535 VOUT.n534 1.13663
R9068 VOUT.n544 VOUT.n543 1.13663
R9069 VOUT.n553 VOUT.n552 1.13663
R9070 VOUT.n562 VOUT.n561 1.13663
R9071 VOUT.n203 VOUT.n202 1.13663
R9072 VOUT.n212 VOUT.n211 1.13663
R9073 VOUT.n221 VOUT.n220 1.13663
R9074 VOUT.n230 VOUT.n229 1.13663
R9075 VOUT.n239 VOUT.n238 1.13663
R9076 VOUT.n248 VOUT.n247 1.13663
R9077 VOUT.n257 VOUT.n256 1.13663
R9078 VOUT.n266 VOUT.n265 1.13663
R9079 VOUT.n275 VOUT.n274 1.13663
R9080 VOUT.n284 VOUT.n283 1.13663
R9081 VOUT.n293 VOUT.n292 1.13663
R9082 VOUT.n302 VOUT.n301 1.13663
R9083 VOUT.n311 VOUT.n310 1.13663
R9084 VOUT.n320 VOUT.n319 1.13663
R9085 VOUT.n329 VOUT.n328 1.13663
R9086 VOUT.n338 VOUT.n337 1.13663
R9087 VOUT.n347 VOUT.n346 1.13663
R9088 VOUT.n356 VOUT.n355 1.13663
R9089 VOUT.n365 VOUT.n364 1.13663
R9090 VOUT.n374 VOUT.n373 1.13663
R9091 VOUT.n15 VOUT.n14 1.13663
R9092 VOUT.n24 VOUT.n23 1.13663
R9093 VOUT.n33 VOUT.n32 1.13663
R9094 VOUT.n42 VOUT.n41 1.13663
R9095 VOUT.n51 VOUT.n50 1.13663
R9096 VOUT.n60 VOUT.n59 1.13663
R9097 VOUT.n69 VOUT.n68 1.13663
R9098 VOUT.n78 VOUT.n77 1.13663
R9099 VOUT.n87 VOUT.n86 1.13663
R9100 VOUT.n96 VOUT.n95 1.13663
R9101 VOUT.n105 VOUT.n104 1.13663
R9102 VOUT.n114 VOUT.n113 1.13663
R9103 VOUT.n123 VOUT.n122 1.13663
R9104 VOUT.n132 VOUT.n131 1.13663
R9105 VOUT.n141 VOUT.n140 1.13663
R9106 VOUT.n150 VOUT.n149 1.13663
R9107 VOUT.n159 VOUT.n158 1.13663
R9108 VOUT.n168 VOUT.n167 1.13663
R9109 VOUT.n177 VOUT.n176 1.13663
R9110 VOUT.n186 VOUT.n185 1.13663
R9111 VOUT.n1691 VOUT.n1690 1.12991
R9112 VOUT.n1682 VOUT.n1681 1.12991
R9113 VOUT.n1673 VOUT.n1672 1.12991
R9114 VOUT.n1664 VOUT.n1663 1.12991
R9115 VOUT.n1655 VOUT.n1654 1.12991
R9116 VOUT.n1646 VOUT.n1645 1.12991
R9117 VOUT.n1637 VOUT.n1636 1.12991
R9118 VOUT.n1628 VOUT.n1627 1.12991
R9119 VOUT.n1619 VOUT.n1618 1.12991
R9120 VOUT.n1610 VOUT.n1609 1.12991
R9121 VOUT.n1601 VOUT.n1600 1.12991
R9122 VOUT.n1592 VOUT.n1591 1.12991
R9123 VOUT.n1583 VOUT.n1582 1.12991
R9124 VOUT.n1574 VOUT.n1573 1.12991
R9125 VOUT.n1565 VOUT.n1564 1.12991
R9126 VOUT.n1556 VOUT.n1555 1.12991
R9127 VOUT.n1547 VOUT.n1546 1.12991
R9128 VOUT.n1538 VOUT.n1537 1.12991
R9129 VOUT.n1529 VOUT.n1528 1.12991
R9130 VOUT.n1520 VOUT.n1519 1.12991
R9131 VOUT.n1511 VOUT.n1510 1.12991
R9132 VOUT.n2455 VOUT.n2454 0.774807
R9133 VOUT.n2455 VOUT.n565 0.501109
R9134 VOUT.n558 VOUT.n557 0.493707
R9135 VOUT.n549 VOUT.n548 0.493707
R9136 VOUT.n540 VOUT.n539 0.493707
R9137 VOUT.n531 VOUT.n530 0.493707
R9138 VOUT.n522 VOUT.n521 0.493707
R9139 VOUT.n513 VOUT.n512 0.493707
R9140 VOUT.n504 VOUT.n503 0.493707
R9141 VOUT.n495 VOUT.n494 0.493707
R9142 VOUT.n486 VOUT.n485 0.493707
R9143 VOUT.n477 VOUT.n476 0.493707
R9144 VOUT.n468 VOUT.n467 0.493707
R9145 VOUT.n459 VOUT.n458 0.493707
R9146 VOUT.n450 VOUT.n449 0.493707
R9147 VOUT.n441 VOUT.n440 0.493707
R9148 VOUT.n432 VOUT.n431 0.493707
R9149 VOUT.n423 VOUT.n422 0.493707
R9150 VOUT.n414 VOUT.n413 0.493707
R9151 VOUT.n405 VOUT.n404 0.493707
R9152 VOUT.n396 VOUT.n395 0.493707
R9153 VOUT.n387 VOUT.n386 0.493707
R9154 VOUT.n379 VOUT.n378 0.493707
R9155 VOUT.n370 VOUT.n369 0.493707
R9156 VOUT.n361 VOUT.n360 0.493707
R9157 VOUT.n352 VOUT.n351 0.493707
R9158 VOUT.n343 VOUT.n342 0.493707
R9159 VOUT.n334 VOUT.n333 0.493707
R9160 VOUT.n325 VOUT.n324 0.493707
R9161 VOUT.n316 VOUT.n315 0.493707
R9162 VOUT.n307 VOUT.n306 0.493707
R9163 VOUT.n298 VOUT.n297 0.493707
R9164 VOUT.n289 VOUT.n288 0.493707
R9165 VOUT.n280 VOUT.n279 0.493707
R9166 VOUT.n271 VOUT.n270 0.493707
R9167 VOUT.n262 VOUT.n261 0.493707
R9168 VOUT.n253 VOUT.n252 0.493707
R9169 VOUT.n244 VOUT.n243 0.493707
R9170 VOUT.n235 VOUT.n234 0.493707
R9171 VOUT.n226 VOUT.n225 0.493707
R9172 VOUT.n217 VOUT.n216 0.493707
R9173 VOUT.n208 VOUT.n207 0.493707
R9174 VOUT.n199 VOUT.n198 0.493707
R9175 VOUT.n191 VOUT.n190 0.493707
R9176 VOUT.n182 VOUT.n181 0.493707
R9177 VOUT.n173 VOUT.n172 0.493707
R9178 VOUT.n164 VOUT.n163 0.493707
R9179 VOUT.n155 VOUT.n154 0.493707
R9180 VOUT.n146 VOUT.n145 0.493707
R9181 VOUT.n137 VOUT.n136 0.493707
R9182 VOUT.n128 VOUT.n127 0.493707
R9183 VOUT.n119 VOUT.n118 0.493707
R9184 VOUT.n110 VOUT.n109 0.493707
R9185 VOUT.n101 VOUT.n100 0.493707
R9186 VOUT.n92 VOUT.n91 0.493707
R9187 VOUT.n83 VOUT.n82 0.493707
R9188 VOUT.n74 VOUT.n73 0.493707
R9189 VOUT.n65 VOUT.n64 0.493707
R9190 VOUT.n56 VOUT.n55 0.493707
R9191 VOUT.n47 VOUT.n46 0.493707
R9192 VOUT.n38 VOUT.n37 0.493707
R9193 VOUT.n29 VOUT.n28 0.493707
R9194 VOUT.n20 VOUT.n19 0.493707
R9195 VOUT.n11 VOUT.n10 0.493707
R9196 VOUT.n3 VOUT.n2 0.493707
R9197 VOUT.n1688 VOUT.n1686 0.394025
R9198 VOUT.n1508 VOUT.n1506 0.394025
R9199 VOUT.n1679 VOUT.n1677 0.394019
R9200 VOUT.n1670 VOUT.n1668 0.394019
R9201 VOUT.n1661 VOUT.n1659 0.394019
R9202 VOUT.n1652 VOUT.n1650 0.394019
R9203 VOUT.n1643 VOUT.n1641 0.394019
R9204 VOUT.n1634 VOUT.n1632 0.394019
R9205 VOUT.n1625 VOUT.n1623 0.394019
R9206 VOUT.n1616 VOUT.n1614 0.394019
R9207 VOUT.n1607 VOUT.n1605 0.394019
R9208 VOUT.n1598 VOUT.n1596 0.394019
R9209 VOUT.n1589 VOUT.n1587 0.394019
R9210 VOUT.n1580 VOUT.n1578 0.394019
R9211 VOUT.n1571 VOUT.n1569 0.394019
R9212 VOUT.n1562 VOUT.n1560 0.394019
R9213 VOUT.n1553 VOUT.n1551 0.394019
R9214 VOUT.n1544 VOUT.n1542 0.394019
R9215 VOUT.n1535 VOUT.n1533 0.394019
R9216 VOUT.n1526 VOUT.n1524 0.394019
R9217 VOUT.n1517 VOUT.n1515 0.394019
R9218 VOUT.n2261 VOUT.n2259 0.37776
R9219 VOUT.n2401 VOUT.n2399 0.37776
R9220 VOUT.n2268 VOUT.n2266 0.377755
R9221 VOUT.n2275 VOUT.n2273 0.377755
R9222 VOUT.n2282 VOUT.n2280 0.377755
R9223 VOUT.n2289 VOUT.n2287 0.377755
R9224 VOUT.n2296 VOUT.n2294 0.377755
R9225 VOUT.n2303 VOUT.n2301 0.377755
R9226 VOUT.n2310 VOUT.n2308 0.377755
R9227 VOUT.n2317 VOUT.n2315 0.377755
R9228 VOUT.n2324 VOUT.n2322 0.377755
R9229 VOUT.n2331 VOUT.n2329 0.377755
R9230 VOUT.n2338 VOUT.n2336 0.377755
R9231 VOUT.n2345 VOUT.n2343 0.377755
R9232 VOUT.n2352 VOUT.n2350 0.377755
R9233 VOUT.n2359 VOUT.n2357 0.377755
R9234 VOUT.n2366 VOUT.n2364 0.377755
R9235 VOUT.n2373 VOUT.n2371 0.377755
R9236 VOUT.n2380 VOUT.n2378 0.377755
R9237 VOUT.n2387 VOUT.n2385 0.377755
R9238 VOUT.n2394 VOUT.n2392 0.377755
R9239 VOUT.n2253 VOUT.n2251 0.366502
R9240 VOUT.n2073 VOUT.n2071 0.366502
R9241 VOUT.n2244 VOUT.n2242 0.366496
R9242 VOUT.n2235 VOUT.n2233 0.366496
R9243 VOUT.n2226 VOUT.n2224 0.366496
R9244 VOUT.n2217 VOUT.n2215 0.366496
R9245 VOUT.n2208 VOUT.n2206 0.366496
R9246 VOUT.n2199 VOUT.n2197 0.366496
R9247 VOUT.n2190 VOUT.n2188 0.366496
R9248 VOUT.n2181 VOUT.n2179 0.366496
R9249 VOUT.n2172 VOUT.n2170 0.366496
R9250 VOUT.n2163 VOUT.n2161 0.366496
R9251 VOUT.n2154 VOUT.n2152 0.366496
R9252 VOUT.n2145 VOUT.n2143 0.366496
R9253 VOUT.n2136 VOUT.n2134 0.366496
R9254 VOUT.n2127 VOUT.n2125 0.366496
R9255 VOUT.n2118 VOUT.n2116 0.366496
R9256 VOUT.n2109 VOUT.n2107 0.366496
R9257 VOUT.n2100 VOUT.n2098 0.366496
R9258 VOUT.n2091 VOUT.n2089 0.366496
R9259 VOUT.n2082 VOUT.n2080 0.366496
R9260 VOUT.n1877 VOUT.n1875 0.360687
R9261 VOUT.n1697 VOUT.n1695 0.360687
R9262 VOUT.n1868 VOUT.n1866 0.360682
R9263 VOUT.n1859 VOUT.n1857 0.360682
R9264 VOUT.n1850 VOUT.n1848 0.360682
R9265 VOUT.n1841 VOUT.n1839 0.360682
R9266 VOUT.n1832 VOUT.n1830 0.360682
R9267 VOUT.n1823 VOUT.n1821 0.360682
R9268 VOUT.n1814 VOUT.n1812 0.360682
R9269 VOUT.n1805 VOUT.n1803 0.360682
R9270 VOUT.n1796 VOUT.n1794 0.360682
R9271 VOUT.n1787 VOUT.n1785 0.360682
R9272 VOUT.n1778 VOUT.n1776 0.360682
R9273 VOUT.n1769 VOUT.n1767 0.360682
R9274 VOUT.n1760 VOUT.n1758 0.360682
R9275 VOUT.n1751 VOUT.n1749 0.360682
R9276 VOUT.n1742 VOUT.n1740 0.360682
R9277 VOUT.n1733 VOUT.n1731 0.360682
R9278 VOUT.n1724 VOUT.n1722 0.360682
R9279 VOUT.n1715 VOUT.n1713 0.360682
R9280 VOUT.n1706 VOUT.n1704 0.360682
R9281 VOUT.n749 VOUT.n747 0.357646
R9282 VOUT.n569 VOUT.n567 0.357646
R9283 VOUT.n2065 VOUT.n2063 0.357646
R9284 VOUT.n1885 VOUT.n1883 0.357646
R9285 VOUT.n740 VOUT.n738 0.35764
R9286 VOUT.n731 VOUT.n729 0.35764
R9287 VOUT.n722 VOUT.n720 0.35764
R9288 VOUT.n713 VOUT.n711 0.35764
R9289 VOUT.n704 VOUT.n702 0.35764
R9290 VOUT.n695 VOUT.n693 0.35764
R9291 VOUT.n686 VOUT.n684 0.35764
R9292 VOUT.n677 VOUT.n675 0.35764
R9293 VOUT.n668 VOUT.n666 0.35764
R9294 VOUT.n659 VOUT.n657 0.35764
R9295 VOUT.n650 VOUT.n648 0.35764
R9296 VOUT.n641 VOUT.n639 0.35764
R9297 VOUT.n632 VOUT.n630 0.35764
R9298 VOUT.n623 VOUT.n621 0.35764
R9299 VOUT.n614 VOUT.n612 0.35764
R9300 VOUT.n605 VOUT.n603 0.35764
R9301 VOUT.n596 VOUT.n594 0.35764
R9302 VOUT.n587 VOUT.n585 0.35764
R9303 VOUT.n578 VOUT.n576 0.35764
R9304 VOUT.n2056 VOUT.n2054 0.35764
R9305 VOUT.n2047 VOUT.n2045 0.35764
R9306 VOUT.n2038 VOUT.n2036 0.35764
R9307 VOUT.n2029 VOUT.n2027 0.35764
R9308 VOUT.n2020 VOUT.n2018 0.35764
R9309 VOUT.n2011 VOUT.n2009 0.35764
R9310 VOUT.n2002 VOUT.n2000 0.35764
R9311 VOUT.n1993 VOUT.n1991 0.35764
R9312 VOUT.n1984 VOUT.n1982 0.35764
R9313 VOUT.n1975 VOUT.n1973 0.35764
R9314 VOUT.n1966 VOUT.n1964 0.35764
R9315 VOUT.n1957 VOUT.n1955 0.35764
R9316 VOUT.n1948 VOUT.n1946 0.35764
R9317 VOUT.n1939 VOUT.n1937 0.35764
R9318 VOUT.n1930 VOUT.n1928 0.35764
R9319 VOUT.n1921 VOUT.n1919 0.35764
R9320 VOUT.n1912 VOUT.n1910 0.35764
R9321 VOUT.n1903 VOUT.n1901 0.35764
R9322 VOUT.n1894 VOUT.n1892 0.35764
R9323 VOUT.n937 VOUT.n935 0.356403
R9324 VOUT.n757 VOUT.n755 0.356403
R9325 VOUT.n928 VOUT.n926 0.356397
R9326 VOUT.n919 VOUT.n917 0.356397
R9327 VOUT.n910 VOUT.n908 0.356397
R9328 VOUT.n901 VOUT.n899 0.356397
R9329 VOUT.n892 VOUT.n890 0.356397
R9330 VOUT.n883 VOUT.n881 0.356397
R9331 VOUT.n874 VOUT.n872 0.356397
R9332 VOUT.n865 VOUT.n863 0.356397
R9333 VOUT.n856 VOUT.n854 0.356397
R9334 VOUT.n847 VOUT.n845 0.356397
R9335 VOUT.n838 VOUT.n836 0.356397
R9336 VOUT.n829 VOUT.n827 0.356397
R9337 VOUT.n820 VOUT.n818 0.356397
R9338 VOUT.n811 VOUT.n809 0.356397
R9339 VOUT.n802 VOUT.n800 0.356397
R9340 VOUT.n793 VOUT.n791 0.356397
R9341 VOUT.n784 VOUT.n782 0.356397
R9342 VOUT.n775 VOUT.n773 0.356397
R9343 VOUT.n766 VOUT.n764 0.356397
R9344 VOUT.n1125 VOUT.n1123 0.353572
R9345 VOUT.n945 VOUT.n943 0.353572
R9346 VOUT.n1116 VOUT.n1114 0.353567
R9347 VOUT.n1107 VOUT.n1105 0.353567
R9348 VOUT.n1098 VOUT.n1096 0.353567
R9349 VOUT.n1089 VOUT.n1087 0.353567
R9350 VOUT.n1080 VOUT.n1078 0.353567
R9351 VOUT.n1071 VOUT.n1069 0.353567
R9352 VOUT.n1062 VOUT.n1060 0.353567
R9353 VOUT.n1053 VOUT.n1051 0.353567
R9354 VOUT.n1044 VOUT.n1042 0.353567
R9355 VOUT.n1035 VOUT.n1033 0.353567
R9356 VOUT.n1026 VOUT.n1024 0.353567
R9357 VOUT.n1017 VOUT.n1015 0.353567
R9358 VOUT.n1008 VOUT.n1006 0.353567
R9359 VOUT.n999 VOUT.n997 0.353567
R9360 VOUT.n990 VOUT.n988 0.353567
R9361 VOUT.n981 VOUT.n979 0.353567
R9362 VOUT.n972 VOUT.n970 0.353567
R9363 VOUT.n963 VOUT.n961 0.353567
R9364 VOUT.n954 VOUT.n952 0.353567
R9365 VOUT.n1313 VOUT.n1311 0.352169
R9366 VOUT.n1133 VOUT.n1131 0.352169
R9367 VOUT.n1304 VOUT.n1302 0.352163
R9368 VOUT.n1295 VOUT.n1293 0.352163
R9369 VOUT.n1286 VOUT.n1284 0.352163
R9370 VOUT.n1277 VOUT.n1275 0.352163
R9371 VOUT.n1268 VOUT.n1266 0.352163
R9372 VOUT.n1259 VOUT.n1257 0.352163
R9373 VOUT.n1250 VOUT.n1248 0.352163
R9374 VOUT.n1241 VOUT.n1239 0.352163
R9375 VOUT.n1232 VOUT.n1230 0.352163
R9376 VOUT.n1223 VOUT.n1221 0.352163
R9377 VOUT.n1214 VOUT.n1212 0.352163
R9378 VOUT.n1205 VOUT.n1203 0.352163
R9379 VOUT.n1196 VOUT.n1194 0.352163
R9380 VOUT.n1187 VOUT.n1185 0.352163
R9381 VOUT.n1178 VOUT.n1176 0.352163
R9382 VOUT.n1169 VOUT.n1167 0.352163
R9383 VOUT.n1160 VOUT.n1158 0.352163
R9384 VOUT.n1151 VOUT.n1149 0.352163
R9385 VOUT.n1142 VOUT.n1140 0.352163
R9386 VOUT.n1501 VOUT.n1499 0.349544
R9387 VOUT.n1321 VOUT.n1319 0.349544
R9388 VOUT.n1492 VOUT.n1490 0.349539
R9389 VOUT.n1483 VOUT.n1481 0.349539
R9390 VOUT.n1474 VOUT.n1472 0.349539
R9391 VOUT.n1465 VOUT.n1463 0.349539
R9392 VOUT.n1456 VOUT.n1454 0.349539
R9393 VOUT.n1447 VOUT.n1445 0.349539
R9394 VOUT.n1438 VOUT.n1436 0.349539
R9395 VOUT.n1429 VOUT.n1427 0.349539
R9396 VOUT.n1420 VOUT.n1418 0.349539
R9397 VOUT.n1411 VOUT.n1409 0.349539
R9398 VOUT.n1402 VOUT.n1400 0.349539
R9399 VOUT.n1393 VOUT.n1391 0.349539
R9400 VOUT.n1384 VOUT.n1382 0.349539
R9401 VOUT.n1375 VOUT.n1373 0.349539
R9402 VOUT.n1366 VOUT.n1364 0.349539
R9403 VOUT.n1357 VOUT.n1355 0.349539
R9404 VOUT.n1348 VOUT.n1346 0.349539
R9405 VOUT.n1339 VOUT.n1337 0.349539
R9406 VOUT.n1330 VOUT.n1328 0.349539
R9407 VOUT.n2446 VOUT.n2445 0.342463
R9408 VOUT.n2450 VOUT.n2449 0.338671
R9409 VOUT.n564 VOUT.n563 0.283561
R9410 VOUT.n2447 VOUT.n2446 0.23963
R9411 VOUT.n2448 VOUT.n2447 0.236913
R9412 VOUT.n2451 VOUT.n2450 0.236913
R9413 VOUT.n2452 VOUT.n2451 0.236913
R9414 VOUT.n2453 VOUT.n2452 0.236913
R9415 VOUT.n2454 VOUT.n2453 0.236913
R9416 VOUT.n745 VOUT.n744 0.236284
R9417 VOUT.n736 VOUT.n735 0.236284
R9418 VOUT.n727 VOUT.n726 0.236284
R9419 VOUT.n718 VOUT.n717 0.236284
R9420 VOUT.n709 VOUT.n708 0.236284
R9421 VOUT.n700 VOUT.n699 0.236284
R9422 VOUT.n691 VOUT.n690 0.236284
R9423 VOUT.n682 VOUT.n681 0.236284
R9424 VOUT.n673 VOUT.n672 0.236284
R9425 VOUT.n664 VOUT.n663 0.236284
R9426 VOUT.n655 VOUT.n654 0.236284
R9427 VOUT.n646 VOUT.n645 0.236284
R9428 VOUT.n637 VOUT.n636 0.236284
R9429 VOUT.n628 VOUT.n627 0.236284
R9430 VOUT.n619 VOUT.n618 0.236284
R9431 VOUT.n610 VOUT.n609 0.236284
R9432 VOUT.n601 VOUT.n600 0.236284
R9433 VOUT.n592 VOUT.n591 0.236284
R9434 VOUT.n583 VOUT.n582 0.236284
R9435 VOUT.n574 VOUT.n573 0.236284
R9436 VOUT.n933 VOUT.n932 0.236284
R9437 VOUT.n924 VOUT.n923 0.236284
R9438 VOUT.n915 VOUT.n914 0.236284
R9439 VOUT.n906 VOUT.n905 0.236284
R9440 VOUT.n897 VOUT.n896 0.236284
R9441 VOUT.n888 VOUT.n887 0.236284
R9442 VOUT.n879 VOUT.n878 0.236284
R9443 VOUT.n870 VOUT.n869 0.236284
R9444 VOUT.n861 VOUT.n860 0.236284
R9445 VOUT.n852 VOUT.n851 0.236284
R9446 VOUT.n843 VOUT.n842 0.236284
R9447 VOUT.n834 VOUT.n833 0.236284
R9448 VOUT.n825 VOUT.n824 0.236284
R9449 VOUT.n816 VOUT.n815 0.236284
R9450 VOUT.n807 VOUT.n806 0.236284
R9451 VOUT.n798 VOUT.n797 0.236284
R9452 VOUT.n789 VOUT.n788 0.236284
R9453 VOUT.n780 VOUT.n779 0.236284
R9454 VOUT.n771 VOUT.n770 0.236284
R9455 VOUT.n762 VOUT.n761 0.236284
R9456 VOUT.n1121 VOUT.n1120 0.236284
R9457 VOUT.n1112 VOUT.n1111 0.236284
R9458 VOUT.n1103 VOUT.n1102 0.236284
R9459 VOUT.n1094 VOUT.n1093 0.236284
R9460 VOUT.n1085 VOUT.n1084 0.236284
R9461 VOUT.n1076 VOUT.n1075 0.236284
R9462 VOUT.n1067 VOUT.n1066 0.236284
R9463 VOUT.n1058 VOUT.n1057 0.236284
R9464 VOUT.n1049 VOUT.n1048 0.236284
R9465 VOUT.n1040 VOUT.n1039 0.236284
R9466 VOUT.n1031 VOUT.n1030 0.236284
R9467 VOUT.n1022 VOUT.n1021 0.236284
R9468 VOUT.n1013 VOUT.n1012 0.236284
R9469 VOUT.n1004 VOUT.n1003 0.236284
R9470 VOUT.n995 VOUT.n994 0.236284
R9471 VOUT.n986 VOUT.n985 0.236284
R9472 VOUT.n977 VOUT.n976 0.236284
R9473 VOUT.n968 VOUT.n967 0.236284
R9474 VOUT.n959 VOUT.n958 0.236284
R9475 VOUT.n950 VOUT.n949 0.236284
R9476 VOUT.n1309 VOUT.n1308 0.236284
R9477 VOUT.n1300 VOUT.n1299 0.236284
R9478 VOUT.n1291 VOUT.n1290 0.236284
R9479 VOUT.n1282 VOUT.n1281 0.236284
R9480 VOUT.n1273 VOUT.n1272 0.236284
R9481 VOUT.n1264 VOUT.n1263 0.236284
R9482 VOUT.n1255 VOUT.n1254 0.236284
R9483 VOUT.n1246 VOUT.n1245 0.236284
R9484 VOUT.n1237 VOUT.n1236 0.236284
R9485 VOUT.n1228 VOUT.n1227 0.236284
R9486 VOUT.n1219 VOUT.n1218 0.236284
R9487 VOUT.n1210 VOUT.n1209 0.236284
R9488 VOUT.n1201 VOUT.n1200 0.236284
R9489 VOUT.n1192 VOUT.n1191 0.236284
R9490 VOUT.n1183 VOUT.n1182 0.236284
R9491 VOUT.n1174 VOUT.n1173 0.236284
R9492 VOUT.n1165 VOUT.n1164 0.236284
R9493 VOUT.n1156 VOUT.n1155 0.236284
R9494 VOUT.n1147 VOUT.n1146 0.236284
R9495 VOUT.n1138 VOUT.n1137 0.236284
R9496 VOUT.n1497 VOUT.n1496 0.236284
R9497 VOUT.n1488 VOUT.n1487 0.236284
R9498 VOUT.n1479 VOUT.n1478 0.236284
R9499 VOUT.n1470 VOUT.n1469 0.236284
R9500 VOUT.n1461 VOUT.n1460 0.236284
R9501 VOUT.n1452 VOUT.n1451 0.236284
R9502 VOUT.n1443 VOUT.n1442 0.236284
R9503 VOUT.n1434 VOUT.n1433 0.236284
R9504 VOUT.n1425 VOUT.n1424 0.236284
R9505 VOUT.n1416 VOUT.n1415 0.236284
R9506 VOUT.n1407 VOUT.n1406 0.236284
R9507 VOUT.n1398 VOUT.n1397 0.236284
R9508 VOUT.n1389 VOUT.n1388 0.236284
R9509 VOUT.n1380 VOUT.n1379 0.236284
R9510 VOUT.n1371 VOUT.n1370 0.236284
R9511 VOUT.n1362 VOUT.n1361 0.236284
R9512 VOUT.n1353 VOUT.n1352 0.236284
R9513 VOUT.n1344 VOUT.n1343 0.236284
R9514 VOUT.n1335 VOUT.n1334 0.236284
R9515 VOUT.n1326 VOUT.n1325 0.236284
R9516 VOUT.n1685 VOUT.n1684 0.236284
R9517 VOUT.n1676 VOUT.n1675 0.236284
R9518 VOUT.n1667 VOUT.n1666 0.236284
R9519 VOUT.n1658 VOUT.n1657 0.236284
R9520 VOUT.n1649 VOUT.n1648 0.236284
R9521 VOUT.n1640 VOUT.n1639 0.236284
R9522 VOUT.n1631 VOUT.n1630 0.236284
R9523 VOUT.n1622 VOUT.n1621 0.236284
R9524 VOUT.n1613 VOUT.n1612 0.236284
R9525 VOUT.n1604 VOUT.n1603 0.236284
R9526 VOUT.n1595 VOUT.n1594 0.236284
R9527 VOUT.n1586 VOUT.n1585 0.236284
R9528 VOUT.n1577 VOUT.n1576 0.236284
R9529 VOUT.n1568 VOUT.n1567 0.236284
R9530 VOUT.n1559 VOUT.n1558 0.236284
R9531 VOUT.n1550 VOUT.n1549 0.236284
R9532 VOUT.n1541 VOUT.n1540 0.236284
R9533 VOUT.n1532 VOUT.n1531 0.236284
R9534 VOUT.n1523 VOUT.n1522 0.236284
R9535 VOUT.n1514 VOUT.n1513 0.236284
R9536 VOUT.n1873 VOUT.n1872 0.236284
R9537 VOUT.n1864 VOUT.n1863 0.236284
R9538 VOUT.n1855 VOUT.n1854 0.236284
R9539 VOUT.n1846 VOUT.n1845 0.236284
R9540 VOUT.n1837 VOUT.n1836 0.236284
R9541 VOUT.n1828 VOUT.n1827 0.236284
R9542 VOUT.n1819 VOUT.n1818 0.236284
R9543 VOUT.n1810 VOUT.n1809 0.236284
R9544 VOUT.n1801 VOUT.n1800 0.236284
R9545 VOUT.n1792 VOUT.n1791 0.236284
R9546 VOUT.n1783 VOUT.n1782 0.236284
R9547 VOUT.n1774 VOUT.n1773 0.236284
R9548 VOUT.n1765 VOUT.n1764 0.236284
R9549 VOUT.n1756 VOUT.n1755 0.236284
R9550 VOUT.n1747 VOUT.n1746 0.236284
R9551 VOUT.n1738 VOUT.n1737 0.236284
R9552 VOUT.n1729 VOUT.n1728 0.236284
R9553 VOUT.n1720 VOUT.n1719 0.236284
R9554 VOUT.n1711 VOUT.n1710 0.236284
R9555 VOUT.n1702 VOUT.n1701 0.236284
R9556 VOUT.n2061 VOUT.n2060 0.236284
R9557 VOUT.n2052 VOUT.n2051 0.236284
R9558 VOUT.n2043 VOUT.n2042 0.236284
R9559 VOUT.n2034 VOUT.n2033 0.236284
R9560 VOUT.n2025 VOUT.n2024 0.236284
R9561 VOUT.n2016 VOUT.n2015 0.236284
R9562 VOUT.n2007 VOUT.n2006 0.236284
R9563 VOUT.n1998 VOUT.n1997 0.236284
R9564 VOUT.n1989 VOUT.n1988 0.236284
R9565 VOUT.n1980 VOUT.n1979 0.236284
R9566 VOUT.n1971 VOUT.n1970 0.236284
R9567 VOUT.n1962 VOUT.n1961 0.236284
R9568 VOUT.n1953 VOUT.n1952 0.236284
R9569 VOUT.n1944 VOUT.n1943 0.236284
R9570 VOUT.n1935 VOUT.n1934 0.236284
R9571 VOUT.n1926 VOUT.n1925 0.236284
R9572 VOUT.n1917 VOUT.n1916 0.236284
R9573 VOUT.n1908 VOUT.n1907 0.236284
R9574 VOUT.n1899 VOUT.n1898 0.236284
R9575 VOUT.n1890 VOUT.n1889 0.236284
R9576 VOUT.n2249 VOUT.n2248 0.236284
R9577 VOUT.n2240 VOUT.n2239 0.236284
R9578 VOUT.n2231 VOUT.n2230 0.236284
R9579 VOUT.n2222 VOUT.n2221 0.236284
R9580 VOUT.n2213 VOUT.n2212 0.236284
R9581 VOUT.n2204 VOUT.n2203 0.236284
R9582 VOUT.n2195 VOUT.n2194 0.236284
R9583 VOUT.n2186 VOUT.n2185 0.236284
R9584 VOUT.n2177 VOUT.n2176 0.236284
R9585 VOUT.n2168 VOUT.n2167 0.236284
R9586 VOUT.n2159 VOUT.n2158 0.236284
R9587 VOUT.n2150 VOUT.n2149 0.236284
R9588 VOUT.n2141 VOUT.n2140 0.236284
R9589 VOUT.n2132 VOUT.n2131 0.236284
R9590 VOUT.n2123 VOUT.n2122 0.236284
R9591 VOUT.n2114 VOUT.n2113 0.236284
R9592 VOUT.n2105 VOUT.n2104 0.236284
R9593 VOUT.n2096 VOUT.n2095 0.236284
R9594 VOUT.n2087 VOUT.n2086 0.236284
R9595 VOUT.n2078 VOUT.n2077 0.236284
R9596 VOUT.n2444 VOUT.n2443 0.236284
R9597 VOUT.n2442 VOUT.n2441 0.236284
R9598 VOUT.n2440 VOUT.n2439 0.236284
R9599 VOUT.n2438 VOUT.n2437 0.236284
R9600 VOUT.n2436 VOUT.n2435 0.236284
R9601 VOUT.n2434 VOUT.n2433 0.236284
R9602 VOUT.n2432 VOUT.n2431 0.236284
R9603 VOUT.n2430 VOUT.n2429 0.236284
R9604 VOUT.n2428 VOUT.n2427 0.236284
R9605 VOUT.n2426 VOUT.n2425 0.236284
R9606 VOUT.n2424 VOUT.n2423 0.236284
R9607 VOUT.n2422 VOUT.n2421 0.236284
R9608 VOUT.n2420 VOUT.n2419 0.236284
R9609 VOUT.n2418 VOUT.n2417 0.236284
R9610 VOUT.n2416 VOUT.n2415 0.236284
R9611 VOUT.n2414 VOUT.n2413 0.236284
R9612 VOUT.n2412 VOUT.n2411 0.236284
R9613 VOUT.n2410 VOUT.n2409 0.236284
R9614 VOUT.n2408 VOUT.n2407 0.236284
R9615 VOUT.n2406 VOUT.n2405 0.236284
R9616 VOUT.n2449 VOUT.n2448 0.231478
R9617 VOUT.n562 VOUT.n554 0.227826
R9618 VOUT.n553 VOUT.n545 0.227826
R9619 VOUT.n544 VOUT.n536 0.227826
R9620 VOUT.n535 VOUT.n527 0.227826
R9621 VOUT.n526 VOUT.n518 0.227826
R9622 VOUT.n517 VOUT.n509 0.227826
R9623 VOUT.n508 VOUT.n500 0.227826
R9624 VOUT.n499 VOUT.n491 0.227826
R9625 VOUT.n490 VOUT.n482 0.227826
R9626 VOUT.n481 VOUT.n473 0.227826
R9627 VOUT.n472 VOUT.n464 0.227826
R9628 VOUT.n463 VOUT.n455 0.227826
R9629 VOUT.n454 VOUT.n446 0.227826
R9630 VOUT.n445 VOUT.n437 0.227826
R9631 VOUT.n436 VOUT.n428 0.227826
R9632 VOUT.n427 VOUT.n419 0.227826
R9633 VOUT.n418 VOUT.n410 0.227826
R9634 VOUT.n409 VOUT.n401 0.227826
R9635 VOUT.n400 VOUT.n392 0.227826
R9636 VOUT.n391 VOUT.n383 0.227826
R9637 VOUT.n374 VOUT.n366 0.227826
R9638 VOUT.n365 VOUT.n357 0.227826
R9639 VOUT.n356 VOUT.n348 0.227826
R9640 VOUT.n347 VOUT.n339 0.227826
R9641 VOUT.n338 VOUT.n330 0.227826
R9642 VOUT.n329 VOUT.n321 0.227826
R9643 VOUT.n320 VOUT.n312 0.227826
R9644 VOUT.n311 VOUT.n303 0.227826
R9645 VOUT.n302 VOUT.n294 0.227826
R9646 VOUT.n293 VOUT.n285 0.227826
R9647 VOUT.n284 VOUT.n276 0.227826
R9648 VOUT.n275 VOUT.n267 0.227826
R9649 VOUT.n266 VOUT.n258 0.227826
R9650 VOUT.n257 VOUT.n249 0.227826
R9651 VOUT.n248 VOUT.n240 0.227826
R9652 VOUT.n239 VOUT.n231 0.227826
R9653 VOUT.n230 VOUT.n222 0.227826
R9654 VOUT.n221 VOUT.n213 0.227826
R9655 VOUT.n212 VOUT.n204 0.227826
R9656 VOUT.n203 VOUT.n195 0.227826
R9657 VOUT.n186 VOUT.n178 0.227826
R9658 VOUT.n177 VOUT.n169 0.227826
R9659 VOUT.n168 VOUT.n160 0.227826
R9660 VOUT.n159 VOUT.n151 0.227826
R9661 VOUT.n150 VOUT.n142 0.227826
R9662 VOUT.n141 VOUT.n133 0.227826
R9663 VOUT.n132 VOUT.n124 0.227826
R9664 VOUT.n123 VOUT.n115 0.227826
R9665 VOUT.n114 VOUT.n106 0.227826
R9666 VOUT.n105 VOUT.n97 0.227826
R9667 VOUT.n96 VOUT.n88 0.227826
R9668 VOUT.n87 VOUT.n79 0.227826
R9669 VOUT.n78 VOUT.n70 0.227826
R9670 VOUT.n69 VOUT.n61 0.227826
R9671 VOUT.n60 VOUT.n52 0.227826
R9672 VOUT.n51 VOUT.n43 0.227826
R9673 VOUT.n42 VOUT.n34 0.227826
R9674 VOUT.n33 VOUT.n25 0.227826
R9675 VOUT.n24 VOUT.n16 0.227826
R9676 VOUT.n15 VOUT.n7 0.227826
R9677 VOUT.n565 VOUT.n564 0.199927
R9678 VOUT.n2454 VOUT.n753 0.103333
R9679 VOUT.n2453 VOUT.n941 0.103333
R9680 VOUT.n2452 VOUT.n1129 0.103333
R9681 VOUT.n2451 VOUT.n1317 0.103333
R9682 VOUT.n2450 VOUT.n1505 0.103333
R9683 VOUT.n2449 VOUT.n1693 0.103333
R9684 VOUT.n2448 VOUT.n1881 0.103333
R9685 VOUT.n2447 VOUT.n2069 0.103333
R9686 VOUT.n2446 VOUT.n2257 0.103333
R9687 VOUT.n564 VOUT.n375 0.0841331
R9688 VOUT.n565 VOUT.n187 0.0841331
R9689 VOUT.n563 VOUT.n562 0.059284
R9690 VOUT.n554 VOUT.n553 0.059284
R9691 VOUT.n545 VOUT.n544 0.059284
R9692 VOUT.n536 VOUT.n535 0.059284
R9693 VOUT.n527 VOUT.n526 0.059284
R9694 VOUT.n518 VOUT.n517 0.059284
R9695 VOUT.n509 VOUT.n508 0.059284
R9696 VOUT.n500 VOUT.n499 0.059284
R9697 VOUT.n491 VOUT.n490 0.059284
R9698 VOUT.n482 VOUT.n481 0.059284
R9699 VOUT.n473 VOUT.n472 0.059284
R9700 VOUT.n464 VOUT.n463 0.059284
R9701 VOUT.n455 VOUT.n454 0.059284
R9702 VOUT.n446 VOUT.n445 0.059284
R9703 VOUT.n437 VOUT.n436 0.059284
R9704 VOUT.n428 VOUT.n427 0.059284
R9705 VOUT.n419 VOUT.n418 0.059284
R9706 VOUT.n410 VOUT.n409 0.059284
R9707 VOUT.n401 VOUT.n400 0.059284
R9708 VOUT.n392 VOUT.n391 0.059284
R9709 VOUT.n375 VOUT.n374 0.059284
R9710 VOUT.n366 VOUT.n365 0.059284
R9711 VOUT.n357 VOUT.n356 0.059284
R9712 VOUT.n348 VOUT.n347 0.059284
R9713 VOUT.n339 VOUT.n338 0.059284
R9714 VOUT.n330 VOUT.n329 0.059284
R9715 VOUT.n321 VOUT.n320 0.059284
R9716 VOUT.n312 VOUT.n311 0.059284
R9717 VOUT.n303 VOUT.n302 0.059284
R9718 VOUT.n294 VOUT.n293 0.059284
R9719 VOUT.n285 VOUT.n284 0.059284
R9720 VOUT.n276 VOUT.n275 0.059284
R9721 VOUT.n267 VOUT.n266 0.059284
R9722 VOUT.n258 VOUT.n257 0.059284
R9723 VOUT.n249 VOUT.n248 0.059284
R9724 VOUT.n240 VOUT.n239 0.059284
R9725 VOUT.n231 VOUT.n230 0.059284
R9726 VOUT.n222 VOUT.n221 0.059284
R9727 VOUT.n213 VOUT.n212 0.059284
R9728 VOUT.n204 VOUT.n203 0.059284
R9729 VOUT.n187 VOUT.n186 0.059284
R9730 VOUT.n178 VOUT.n177 0.059284
R9731 VOUT.n169 VOUT.n168 0.059284
R9732 VOUT.n160 VOUT.n159 0.059284
R9733 VOUT.n151 VOUT.n150 0.059284
R9734 VOUT.n142 VOUT.n141 0.059284
R9735 VOUT.n133 VOUT.n132 0.059284
R9736 VOUT.n124 VOUT.n123 0.059284
R9737 VOUT.n115 VOUT.n114 0.059284
R9738 VOUT.n106 VOUT.n105 0.059284
R9739 VOUT.n97 VOUT.n96 0.059284
R9740 VOUT.n88 VOUT.n87 0.059284
R9741 VOUT.n79 VOUT.n78 0.059284
R9742 VOUT.n70 VOUT.n69 0.059284
R9743 VOUT.n61 VOUT.n60 0.059284
R9744 VOUT.n52 VOUT.n51 0.059284
R9745 VOUT.n43 VOUT.n42 0.059284
R9746 VOUT.n34 VOUT.n33 0.059284
R9747 VOUT.n25 VOUT.n24 0.059284
R9748 VOUT.n16 VOUT.n15 0.059284
R9749 VOUT.n753 VOUT.n745 0.0527417
R9750 VOUT.n744 VOUT.n736 0.0527417
R9751 VOUT.n735 VOUT.n727 0.0527417
R9752 VOUT.n726 VOUT.n718 0.0527417
R9753 VOUT.n717 VOUT.n709 0.0527417
R9754 VOUT.n708 VOUT.n700 0.0527417
R9755 VOUT.n699 VOUT.n691 0.0527417
R9756 VOUT.n690 VOUT.n682 0.0527417
R9757 VOUT.n681 VOUT.n673 0.0527417
R9758 VOUT.n672 VOUT.n664 0.0527417
R9759 VOUT.n663 VOUT.n655 0.0527417
R9760 VOUT.n654 VOUT.n646 0.0527417
R9761 VOUT.n645 VOUT.n637 0.0527417
R9762 VOUT.n636 VOUT.n628 0.0527417
R9763 VOUT.n627 VOUT.n619 0.0527417
R9764 VOUT.n618 VOUT.n610 0.0527417
R9765 VOUT.n609 VOUT.n601 0.0527417
R9766 VOUT.n600 VOUT.n592 0.0527417
R9767 VOUT.n591 VOUT.n583 0.0527417
R9768 VOUT.n582 VOUT.n574 0.0527417
R9769 VOUT.n941 VOUT.n933 0.0527417
R9770 VOUT.n932 VOUT.n924 0.0527417
R9771 VOUT.n923 VOUT.n915 0.0527417
R9772 VOUT.n914 VOUT.n906 0.0527417
R9773 VOUT.n905 VOUT.n897 0.0527417
R9774 VOUT.n896 VOUT.n888 0.0527417
R9775 VOUT.n887 VOUT.n879 0.0527417
R9776 VOUT.n878 VOUT.n870 0.0527417
R9777 VOUT.n869 VOUT.n861 0.0527417
R9778 VOUT.n860 VOUT.n852 0.0527417
R9779 VOUT.n851 VOUT.n843 0.0527417
R9780 VOUT.n842 VOUT.n834 0.0527417
R9781 VOUT.n833 VOUT.n825 0.0527417
R9782 VOUT.n824 VOUT.n816 0.0527417
R9783 VOUT.n815 VOUT.n807 0.0527417
R9784 VOUT.n806 VOUT.n798 0.0527417
R9785 VOUT.n797 VOUT.n789 0.0527417
R9786 VOUT.n788 VOUT.n780 0.0527417
R9787 VOUT.n779 VOUT.n771 0.0527417
R9788 VOUT.n770 VOUT.n762 0.0527417
R9789 VOUT.n1129 VOUT.n1121 0.0527417
R9790 VOUT.n1120 VOUT.n1112 0.0527417
R9791 VOUT.n1111 VOUT.n1103 0.0527417
R9792 VOUT.n1102 VOUT.n1094 0.0527417
R9793 VOUT.n1093 VOUT.n1085 0.0527417
R9794 VOUT.n1084 VOUT.n1076 0.0527417
R9795 VOUT.n1075 VOUT.n1067 0.0527417
R9796 VOUT.n1066 VOUT.n1058 0.0527417
R9797 VOUT.n1057 VOUT.n1049 0.0527417
R9798 VOUT.n1048 VOUT.n1040 0.0527417
R9799 VOUT.n1039 VOUT.n1031 0.0527417
R9800 VOUT.n1030 VOUT.n1022 0.0527417
R9801 VOUT.n1021 VOUT.n1013 0.0527417
R9802 VOUT.n1012 VOUT.n1004 0.0527417
R9803 VOUT.n1003 VOUT.n995 0.0527417
R9804 VOUT.n994 VOUT.n986 0.0527417
R9805 VOUT.n985 VOUT.n977 0.0527417
R9806 VOUT.n976 VOUT.n968 0.0527417
R9807 VOUT.n967 VOUT.n959 0.0527417
R9808 VOUT.n958 VOUT.n950 0.0527417
R9809 VOUT.n1317 VOUT.n1309 0.0527417
R9810 VOUT.n1308 VOUT.n1300 0.0527417
R9811 VOUT.n1299 VOUT.n1291 0.0527417
R9812 VOUT.n1290 VOUT.n1282 0.0527417
R9813 VOUT.n1281 VOUT.n1273 0.0527417
R9814 VOUT.n1272 VOUT.n1264 0.0527417
R9815 VOUT.n1263 VOUT.n1255 0.0527417
R9816 VOUT.n1254 VOUT.n1246 0.0527417
R9817 VOUT.n1245 VOUT.n1237 0.0527417
R9818 VOUT.n1236 VOUT.n1228 0.0527417
R9819 VOUT.n1227 VOUT.n1219 0.0527417
R9820 VOUT.n1218 VOUT.n1210 0.0527417
R9821 VOUT.n1209 VOUT.n1201 0.0527417
R9822 VOUT.n1200 VOUT.n1192 0.0527417
R9823 VOUT.n1191 VOUT.n1183 0.0527417
R9824 VOUT.n1182 VOUT.n1174 0.0527417
R9825 VOUT.n1173 VOUT.n1165 0.0527417
R9826 VOUT.n1164 VOUT.n1156 0.0527417
R9827 VOUT.n1155 VOUT.n1147 0.0527417
R9828 VOUT.n1146 VOUT.n1138 0.0527417
R9829 VOUT.n1505 VOUT.n1497 0.0527417
R9830 VOUT.n1496 VOUT.n1488 0.0527417
R9831 VOUT.n1487 VOUT.n1479 0.0527417
R9832 VOUT.n1478 VOUT.n1470 0.0527417
R9833 VOUT.n1469 VOUT.n1461 0.0527417
R9834 VOUT.n1460 VOUT.n1452 0.0527417
R9835 VOUT.n1451 VOUT.n1443 0.0527417
R9836 VOUT.n1442 VOUT.n1434 0.0527417
R9837 VOUT.n1433 VOUT.n1425 0.0527417
R9838 VOUT.n1424 VOUT.n1416 0.0527417
R9839 VOUT.n1415 VOUT.n1407 0.0527417
R9840 VOUT.n1406 VOUT.n1398 0.0527417
R9841 VOUT.n1397 VOUT.n1389 0.0527417
R9842 VOUT.n1388 VOUT.n1380 0.0527417
R9843 VOUT.n1379 VOUT.n1371 0.0527417
R9844 VOUT.n1370 VOUT.n1362 0.0527417
R9845 VOUT.n1361 VOUT.n1353 0.0527417
R9846 VOUT.n1352 VOUT.n1344 0.0527417
R9847 VOUT.n1343 VOUT.n1335 0.0527417
R9848 VOUT.n1334 VOUT.n1326 0.0527417
R9849 VOUT.n1693 VOUT.n1685 0.0527417
R9850 VOUT.n1684 VOUT.n1676 0.0527417
R9851 VOUT.n1675 VOUT.n1667 0.0527417
R9852 VOUT.n1666 VOUT.n1658 0.0527417
R9853 VOUT.n1657 VOUT.n1649 0.0527417
R9854 VOUT.n1648 VOUT.n1640 0.0527417
R9855 VOUT.n1639 VOUT.n1631 0.0527417
R9856 VOUT.n1630 VOUT.n1622 0.0527417
R9857 VOUT.n1621 VOUT.n1613 0.0527417
R9858 VOUT.n1612 VOUT.n1604 0.0527417
R9859 VOUT.n1603 VOUT.n1595 0.0527417
R9860 VOUT.n1594 VOUT.n1586 0.0527417
R9861 VOUT.n1585 VOUT.n1577 0.0527417
R9862 VOUT.n1576 VOUT.n1568 0.0527417
R9863 VOUT.n1567 VOUT.n1559 0.0527417
R9864 VOUT.n1558 VOUT.n1550 0.0527417
R9865 VOUT.n1549 VOUT.n1541 0.0527417
R9866 VOUT.n1540 VOUT.n1532 0.0527417
R9867 VOUT.n1531 VOUT.n1523 0.0527417
R9868 VOUT.n1522 VOUT.n1514 0.0527417
R9869 VOUT.n1881 VOUT.n1873 0.0527417
R9870 VOUT.n1872 VOUT.n1864 0.0527417
R9871 VOUT.n1863 VOUT.n1855 0.0527417
R9872 VOUT.n1854 VOUT.n1846 0.0527417
R9873 VOUT.n1845 VOUT.n1837 0.0527417
R9874 VOUT.n1836 VOUT.n1828 0.0527417
R9875 VOUT.n1827 VOUT.n1819 0.0527417
R9876 VOUT.n1818 VOUT.n1810 0.0527417
R9877 VOUT.n1809 VOUT.n1801 0.0527417
R9878 VOUT.n1800 VOUT.n1792 0.0527417
R9879 VOUT.n1791 VOUT.n1783 0.0527417
R9880 VOUT.n1782 VOUT.n1774 0.0527417
R9881 VOUT.n1773 VOUT.n1765 0.0527417
R9882 VOUT.n1764 VOUT.n1756 0.0527417
R9883 VOUT.n1755 VOUT.n1747 0.0527417
R9884 VOUT.n1746 VOUT.n1738 0.0527417
R9885 VOUT.n1737 VOUT.n1729 0.0527417
R9886 VOUT.n1728 VOUT.n1720 0.0527417
R9887 VOUT.n1719 VOUT.n1711 0.0527417
R9888 VOUT.n1710 VOUT.n1702 0.0527417
R9889 VOUT.n2069 VOUT.n2061 0.0527417
R9890 VOUT.n2060 VOUT.n2052 0.0527417
R9891 VOUT.n2051 VOUT.n2043 0.0527417
R9892 VOUT.n2042 VOUT.n2034 0.0527417
R9893 VOUT.n2033 VOUT.n2025 0.0527417
R9894 VOUT.n2024 VOUT.n2016 0.0527417
R9895 VOUT.n2015 VOUT.n2007 0.0527417
R9896 VOUT.n2006 VOUT.n1998 0.0527417
R9897 VOUT.n1997 VOUT.n1989 0.0527417
R9898 VOUT.n1988 VOUT.n1980 0.0527417
R9899 VOUT.n1979 VOUT.n1971 0.0527417
R9900 VOUT.n1970 VOUT.n1962 0.0527417
R9901 VOUT.n1961 VOUT.n1953 0.0527417
R9902 VOUT.n1952 VOUT.n1944 0.0527417
R9903 VOUT.n1943 VOUT.n1935 0.0527417
R9904 VOUT.n1934 VOUT.n1926 0.0527417
R9905 VOUT.n1925 VOUT.n1917 0.0527417
R9906 VOUT.n1916 VOUT.n1908 0.0527417
R9907 VOUT.n1907 VOUT.n1899 0.0527417
R9908 VOUT.n1898 VOUT.n1890 0.0527417
R9909 VOUT.n2257 VOUT.n2249 0.0527417
R9910 VOUT.n2248 VOUT.n2240 0.0527417
R9911 VOUT.n2239 VOUT.n2231 0.0527417
R9912 VOUT.n2230 VOUT.n2222 0.0527417
R9913 VOUT.n2221 VOUT.n2213 0.0527417
R9914 VOUT.n2212 VOUT.n2204 0.0527417
R9915 VOUT.n2203 VOUT.n2195 0.0527417
R9916 VOUT.n2194 VOUT.n2186 0.0527417
R9917 VOUT.n2185 VOUT.n2177 0.0527417
R9918 VOUT.n2176 VOUT.n2168 0.0527417
R9919 VOUT.n2167 VOUT.n2159 0.0527417
R9920 VOUT.n2158 VOUT.n2150 0.0527417
R9921 VOUT.n2149 VOUT.n2141 0.0527417
R9922 VOUT.n2140 VOUT.n2132 0.0527417
R9923 VOUT.n2131 VOUT.n2123 0.0527417
R9924 VOUT.n2122 VOUT.n2114 0.0527417
R9925 VOUT.n2113 VOUT.n2105 0.0527417
R9926 VOUT.n2104 VOUT.n2096 0.0527417
R9927 VOUT.n2095 VOUT.n2087 0.0527417
R9928 VOUT.n2086 VOUT.n2078 0.0527417
R9929 VOUT.n2445 VOUT.n2444 0.0527417
R9930 VOUT.n2443 VOUT.n2442 0.0527417
R9931 VOUT.n2441 VOUT.n2440 0.0527417
R9932 VOUT.n2439 VOUT.n2438 0.0527417
R9933 VOUT.n2437 VOUT.n2436 0.0527417
R9934 VOUT.n2435 VOUT.n2434 0.0527417
R9935 VOUT.n2433 VOUT.n2432 0.0527417
R9936 VOUT.n2431 VOUT.n2430 0.0527417
R9937 VOUT.n2429 VOUT.n2428 0.0527417
R9938 VOUT.n2427 VOUT.n2426 0.0527417
R9939 VOUT.n2425 VOUT.n2424 0.0527417
R9940 VOUT.n2423 VOUT.n2422 0.0527417
R9941 VOUT.n2421 VOUT.n2420 0.0527417
R9942 VOUT.n2419 VOUT.n2418 0.0527417
R9943 VOUT.n2417 VOUT.n2416 0.0527417
R9944 VOUT.n2415 VOUT.n2414 0.0527417
R9945 VOUT.n2413 VOUT.n2412 0.0527417
R9946 VOUT.n2411 VOUT.n2410 0.0527417
R9947 VOUT.n2409 VOUT.n2408 0.0527417
R9948 VOUT.n2407 VOUT.n2406 0.0527417
R9949 VOUT VOUT.n2455 0.0304363
R9950 VOUT.n558 VOUT.n555 0.0278438
R9951 VOUT.n549 VOUT.n546 0.0278438
R9952 VOUT.n540 VOUT.n537 0.0278438
R9953 VOUT.n531 VOUT.n528 0.0278438
R9954 VOUT.n522 VOUT.n519 0.0278438
R9955 VOUT.n513 VOUT.n510 0.0278438
R9956 VOUT.n504 VOUT.n501 0.0278438
R9957 VOUT.n495 VOUT.n492 0.0278438
R9958 VOUT.n486 VOUT.n483 0.0278438
R9959 VOUT.n477 VOUT.n474 0.0278438
R9960 VOUT.n468 VOUT.n465 0.0278438
R9961 VOUT.n459 VOUT.n456 0.0278438
R9962 VOUT.n450 VOUT.n447 0.0278438
R9963 VOUT.n441 VOUT.n438 0.0278438
R9964 VOUT.n432 VOUT.n429 0.0278438
R9965 VOUT.n423 VOUT.n420 0.0278438
R9966 VOUT.n414 VOUT.n411 0.0278438
R9967 VOUT.n405 VOUT.n402 0.0278438
R9968 VOUT.n396 VOUT.n393 0.0278438
R9969 VOUT.n387 VOUT.n384 0.0278438
R9970 VOUT.n379 VOUT.n376 0.0278438
R9971 VOUT.n370 VOUT.n367 0.0278438
R9972 VOUT.n361 VOUT.n358 0.0278438
R9973 VOUT.n352 VOUT.n349 0.0278438
R9974 VOUT.n343 VOUT.n340 0.0278438
R9975 VOUT.n334 VOUT.n331 0.0278438
R9976 VOUT.n325 VOUT.n322 0.0278438
R9977 VOUT.n316 VOUT.n313 0.0278438
R9978 VOUT.n307 VOUT.n304 0.0278438
R9979 VOUT.n298 VOUT.n295 0.0278438
R9980 VOUT.n289 VOUT.n286 0.0278438
R9981 VOUT.n280 VOUT.n277 0.0278438
R9982 VOUT.n271 VOUT.n268 0.0278438
R9983 VOUT.n262 VOUT.n259 0.0278438
R9984 VOUT.n253 VOUT.n250 0.0278438
R9985 VOUT.n244 VOUT.n241 0.0278438
R9986 VOUT.n235 VOUT.n232 0.0278438
R9987 VOUT.n226 VOUT.n223 0.0278438
R9988 VOUT.n217 VOUT.n214 0.0278438
R9989 VOUT.n208 VOUT.n205 0.0278438
R9990 VOUT.n199 VOUT.n196 0.0278438
R9991 VOUT.n191 VOUT.n188 0.0278438
R9992 VOUT.n182 VOUT.n179 0.0278438
R9993 VOUT.n173 VOUT.n170 0.0278438
R9994 VOUT.n164 VOUT.n161 0.0278438
R9995 VOUT.n155 VOUT.n152 0.0278438
R9996 VOUT.n146 VOUT.n143 0.0278438
R9997 VOUT.n137 VOUT.n134 0.0278438
R9998 VOUT.n128 VOUT.n125 0.0278438
R9999 VOUT.n119 VOUT.n116 0.0278438
R10000 VOUT.n110 VOUT.n107 0.0278438
R10001 VOUT.n101 VOUT.n98 0.0278438
R10002 VOUT.n92 VOUT.n89 0.0278438
R10003 VOUT.n83 VOUT.n80 0.0278438
R10004 VOUT.n74 VOUT.n71 0.0278438
R10005 VOUT.n65 VOUT.n62 0.0278438
R10006 VOUT.n56 VOUT.n53 0.0278438
R10007 VOUT.n47 VOUT.n44 0.0278438
R10008 VOUT.n38 VOUT.n35 0.0278438
R10009 VOUT.n29 VOUT.n26 0.0278438
R10010 VOUT.n20 VOUT.n17 0.0278438
R10011 VOUT.n11 VOUT.n8 0.0278438
R10012 VOUT.n3 VOUT.n0 0.0278438
R10013 VOUT.n749 VOUT.n748 0.0219844
R10014 VOUT.n740 VOUT.n739 0.0219844
R10015 VOUT.n731 VOUT.n730 0.0219844
R10016 VOUT.n722 VOUT.n721 0.0219844
R10017 VOUT.n713 VOUT.n712 0.0219844
R10018 VOUT.n704 VOUT.n703 0.0219844
R10019 VOUT.n695 VOUT.n694 0.0219844
R10020 VOUT.n686 VOUT.n685 0.0219844
R10021 VOUT.n677 VOUT.n676 0.0219844
R10022 VOUT.n668 VOUT.n667 0.0219844
R10023 VOUT.n659 VOUT.n658 0.0219844
R10024 VOUT.n650 VOUT.n649 0.0219844
R10025 VOUT.n641 VOUT.n640 0.0219844
R10026 VOUT.n632 VOUT.n631 0.0219844
R10027 VOUT.n623 VOUT.n622 0.0219844
R10028 VOUT.n614 VOUT.n613 0.0219844
R10029 VOUT.n605 VOUT.n604 0.0219844
R10030 VOUT.n596 VOUT.n595 0.0219844
R10031 VOUT.n587 VOUT.n586 0.0219844
R10032 VOUT.n578 VOUT.n577 0.0219844
R10033 VOUT.n569 VOUT.n568 0.0219844
R10034 VOUT.n937 VOUT.n936 0.0219844
R10035 VOUT.n928 VOUT.n927 0.0219844
R10036 VOUT.n919 VOUT.n918 0.0219844
R10037 VOUT.n910 VOUT.n909 0.0219844
R10038 VOUT.n901 VOUT.n900 0.0219844
R10039 VOUT.n892 VOUT.n891 0.0219844
R10040 VOUT.n883 VOUT.n882 0.0219844
R10041 VOUT.n874 VOUT.n873 0.0219844
R10042 VOUT.n865 VOUT.n864 0.0219844
R10043 VOUT.n856 VOUT.n855 0.0219844
R10044 VOUT.n847 VOUT.n846 0.0219844
R10045 VOUT.n838 VOUT.n837 0.0219844
R10046 VOUT.n829 VOUT.n828 0.0219844
R10047 VOUT.n820 VOUT.n819 0.0219844
R10048 VOUT.n811 VOUT.n810 0.0219844
R10049 VOUT.n802 VOUT.n801 0.0219844
R10050 VOUT.n793 VOUT.n792 0.0219844
R10051 VOUT.n784 VOUT.n783 0.0219844
R10052 VOUT.n775 VOUT.n774 0.0219844
R10053 VOUT.n766 VOUT.n765 0.0219844
R10054 VOUT.n757 VOUT.n756 0.0219844
R10055 VOUT.n1125 VOUT.n1124 0.0219844
R10056 VOUT.n1116 VOUT.n1115 0.0219844
R10057 VOUT.n1107 VOUT.n1106 0.0219844
R10058 VOUT.n1098 VOUT.n1097 0.0219844
R10059 VOUT.n1089 VOUT.n1088 0.0219844
R10060 VOUT.n1080 VOUT.n1079 0.0219844
R10061 VOUT.n1071 VOUT.n1070 0.0219844
R10062 VOUT.n1062 VOUT.n1061 0.0219844
R10063 VOUT.n1053 VOUT.n1052 0.0219844
R10064 VOUT.n1044 VOUT.n1043 0.0219844
R10065 VOUT.n1035 VOUT.n1034 0.0219844
R10066 VOUT.n1026 VOUT.n1025 0.0219844
R10067 VOUT.n1017 VOUT.n1016 0.0219844
R10068 VOUT.n1008 VOUT.n1007 0.0219844
R10069 VOUT.n999 VOUT.n998 0.0219844
R10070 VOUT.n990 VOUT.n989 0.0219844
R10071 VOUT.n981 VOUT.n980 0.0219844
R10072 VOUT.n972 VOUT.n971 0.0219844
R10073 VOUT.n963 VOUT.n962 0.0219844
R10074 VOUT.n954 VOUT.n953 0.0219844
R10075 VOUT.n945 VOUT.n944 0.0219844
R10076 VOUT.n1313 VOUT.n1312 0.0219844
R10077 VOUT.n1304 VOUT.n1303 0.0219844
R10078 VOUT.n1295 VOUT.n1294 0.0219844
R10079 VOUT.n1286 VOUT.n1285 0.0219844
R10080 VOUT.n1277 VOUT.n1276 0.0219844
R10081 VOUT.n1268 VOUT.n1267 0.0219844
R10082 VOUT.n1259 VOUT.n1258 0.0219844
R10083 VOUT.n1250 VOUT.n1249 0.0219844
R10084 VOUT.n1241 VOUT.n1240 0.0219844
R10085 VOUT.n1232 VOUT.n1231 0.0219844
R10086 VOUT.n1223 VOUT.n1222 0.0219844
R10087 VOUT.n1214 VOUT.n1213 0.0219844
R10088 VOUT.n1205 VOUT.n1204 0.0219844
R10089 VOUT.n1196 VOUT.n1195 0.0219844
R10090 VOUT.n1187 VOUT.n1186 0.0219844
R10091 VOUT.n1178 VOUT.n1177 0.0219844
R10092 VOUT.n1169 VOUT.n1168 0.0219844
R10093 VOUT.n1160 VOUT.n1159 0.0219844
R10094 VOUT.n1151 VOUT.n1150 0.0219844
R10095 VOUT.n1142 VOUT.n1141 0.0219844
R10096 VOUT.n1133 VOUT.n1132 0.0219844
R10097 VOUT.n1501 VOUT.n1500 0.0219844
R10098 VOUT.n1492 VOUT.n1491 0.0219844
R10099 VOUT.n1483 VOUT.n1482 0.0219844
R10100 VOUT.n1474 VOUT.n1473 0.0219844
R10101 VOUT.n1465 VOUT.n1464 0.0219844
R10102 VOUT.n1456 VOUT.n1455 0.0219844
R10103 VOUT.n1447 VOUT.n1446 0.0219844
R10104 VOUT.n1438 VOUT.n1437 0.0219844
R10105 VOUT.n1429 VOUT.n1428 0.0219844
R10106 VOUT.n1420 VOUT.n1419 0.0219844
R10107 VOUT.n1411 VOUT.n1410 0.0219844
R10108 VOUT.n1402 VOUT.n1401 0.0219844
R10109 VOUT.n1393 VOUT.n1392 0.0219844
R10110 VOUT.n1384 VOUT.n1383 0.0219844
R10111 VOUT.n1375 VOUT.n1374 0.0219844
R10112 VOUT.n1366 VOUT.n1365 0.0219844
R10113 VOUT.n1357 VOUT.n1356 0.0219844
R10114 VOUT.n1348 VOUT.n1347 0.0219844
R10115 VOUT.n1339 VOUT.n1338 0.0219844
R10116 VOUT.n1330 VOUT.n1329 0.0219844
R10117 VOUT.n1321 VOUT.n1320 0.0219844
R10118 VOUT.n1688 VOUT.n1687 0.0219844
R10119 VOUT.n1679 VOUT.n1678 0.0219844
R10120 VOUT.n1670 VOUT.n1669 0.0219844
R10121 VOUT.n1661 VOUT.n1660 0.0219844
R10122 VOUT.n1652 VOUT.n1651 0.0219844
R10123 VOUT.n1643 VOUT.n1642 0.0219844
R10124 VOUT.n1634 VOUT.n1633 0.0219844
R10125 VOUT.n1625 VOUT.n1624 0.0219844
R10126 VOUT.n1616 VOUT.n1615 0.0219844
R10127 VOUT.n1607 VOUT.n1606 0.0219844
R10128 VOUT.n1598 VOUT.n1597 0.0219844
R10129 VOUT.n1589 VOUT.n1588 0.0219844
R10130 VOUT.n1580 VOUT.n1579 0.0219844
R10131 VOUT.n1571 VOUT.n1570 0.0219844
R10132 VOUT.n1562 VOUT.n1561 0.0219844
R10133 VOUT.n1553 VOUT.n1552 0.0219844
R10134 VOUT.n1544 VOUT.n1543 0.0219844
R10135 VOUT.n1535 VOUT.n1534 0.0219844
R10136 VOUT.n1526 VOUT.n1525 0.0219844
R10137 VOUT.n1517 VOUT.n1516 0.0219844
R10138 VOUT.n1508 VOUT.n1507 0.0219844
R10139 VOUT.n1877 VOUT.n1876 0.0219844
R10140 VOUT.n1868 VOUT.n1867 0.0219844
R10141 VOUT.n1859 VOUT.n1858 0.0219844
R10142 VOUT.n1850 VOUT.n1849 0.0219844
R10143 VOUT.n1841 VOUT.n1840 0.0219844
R10144 VOUT.n1832 VOUT.n1831 0.0219844
R10145 VOUT.n1823 VOUT.n1822 0.0219844
R10146 VOUT.n1814 VOUT.n1813 0.0219844
R10147 VOUT.n1805 VOUT.n1804 0.0219844
R10148 VOUT.n1796 VOUT.n1795 0.0219844
R10149 VOUT.n1787 VOUT.n1786 0.0219844
R10150 VOUT.n1778 VOUT.n1777 0.0219844
R10151 VOUT.n1769 VOUT.n1768 0.0219844
R10152 VOUT.n1760 VOUT.n1759 0.0219844
R10153 VOUT.n1751 VOUT.n1750 0.0219844
R10154 VOUT.n1742 VOUT.n1741 0.0219844
R10155 VOUT.n1733 VOUT.n1732 0.0219844
R10156 VOUT.n1724 VOUT.n1723 0.0219844
R10157 VOUT.n1715 VOUT.n1714 0.0219844
R10158 VOUT.n1706 VOUT.n1705 0.0219844
R10159 VOUT.n1697 VOUT.n1696 0.0219844
R10160 VOUT.n2065 VOUT.n2064 0.0219844
R10161 VOUT.n2056 VOUT.n2055 0.0219844
R10162 VOUT.n2047 VOUT.n2046 0.0219844
R10163 VOUT.n2038 VOUT.n2037 0.0219844
R10164 VOUT.n2029 VOUT.n2028 0.0219844
R10165 VOUT.n2020 VOUT.n2019 0.0219844
R10166 VOUT.n2011 VOUT.n2010 0.0219844
R10167 VOUT.n2002 VOUT.n2001 0.0219844
R10168 VOUT.n1993 VOUT.n1992 0.0219844
R10169 VOUT.n1984 VOUT.n1983 0.0219844
R10170 VOUT.n1975 VOUT.n1974 0.0219844
R10171 VOUT.n1966 VOUT.n1965 0.0219844
R10172 VOUT.n1957 VOUT.n1956 0.0219844
R10173 VOUT.n1948 VOUT.n1947 0.0219844
R10174 VOUT.n1939 VOUT.n1938 0.0219844
R10175 VOUT.n1930 VOUT.n1929 0.0219844
R10176 VOUT.n1921 VOUT.n1920 0.0219844
R10177 VOUT.n1912 VOUT.n1911 0.0219844
R10178 VOUT.n1903 VOUT.n1902 0.0219844
R10179 VOUT.n1894 VOUT.n1893 0.0219844
R10180 VOUT.n1885 VOUT.n1884 0.0219844
R10181 VOUT.n2253 VOUT.n2252 0.0219844
R10182 VOUT.n2244 VOUT.n2243 0.0219844
R10183 VOUT.n2235 VOUT.n2234 0.0219844
R10184 VOUT.n2226 VOUT.n2225 0.0219844
R10185 VOUT.n2217 VOUT.n2216 0.0219844
R10186 VOUT.n2208 VOUT.n2207 0.0219844
R10187 VOUT.n2199 VOUT.n2198 0.0219844
R10188 VOUT.n2190 VOUT.n2189 0.0219844
R10189 VOUT.n2181 VOUT.n2180 0.0219844
R10190 VOUT.n2172 VOUT.n2171 0.0219844
R10191 VOUT.n2163 VOUT.n2162 0.0219844
R10192 VOUT.n2154 VOUT.n2153 0.0219844
R10193 VOUT.n2145 VOUT.n2144 0.0219844
R10194 VOUT.n2136 VOUT.n2135 0.0219844
R10195 VOUT.n2127 VOUT.n2126 0.0219844
R10196 VOUT.n2118 VOUT.n2117 0.0219844
R10197 VOUT.n2109 VOUT.n2108 0.0219844
R10198 VOUT.n2100 VOUT.n2099 0.0219844
R10199 VOUT.n2091 VOUT.n2090 0.0219844
R10200 VOUT.n2082 VOUT.n2081 0.0219844
R10201 VOUT.n2073 VOUT.n2072 0.0219844
R10202 VOUT.n2261 VOUT.n2260 0.0219844
R10203 VOUT.n2268 VOUT.n2267 0.0219844
R10204 VOUT.n2275 VOUT.n2274 0.0219844
R10205 VOUT.n2282 VOUT.n2281 0.0219844
R10206 VOUT.n2289 VOUT.n2288 0.0219844
R10207 VOUT.n2296 VOUT.n2295 0.0219844
R10208 VOUT.n2303 VOUT.n2302 0.0219844
R10209 VOUT.n2310 VOUT.n2309 0.0219844
R10210 VOUT.n2317 VOUT.n2316 0.0219844
R10211 VOUT.n2324 VOUT.n2323 0.0219844
R10212 VOUT.n2331 VOUT.n2330 0.0219844
R10213 VOUT.n2338 VOUT.n2337 0.0219844
R10214 VOUT.n2345 VOUT.n2344 0.0219844
R10215 VOUT.n2352 VOUT.n2351 0.0219844
R10216 VOUT.n2359 VOUT.n2358 0.0219844
R10217 VOUT.n2366 VOUT.n2365 0.0219844
R10218 VOUT.n2373 VOUT.n2372 0.0219844
R10219 VOUT.n2380 VOUT.n2379 0.0219844
R10220 VOUT.n2387 VOUT.n2386 0.0219844
R10221 VOUT.n2394 VOUT.n2393 0.0219844
R10222 VOUT.n2401 VOUT.n2400 0.0219844
R10223 VOUT.n752 VOUT.n749 0.0174092
R10224 VOUT.n743 VOUT.n740 0.0174092
R10225 VOUT.n734 VOUT.n731 0.0174092
R10226 VOUT.n725 VOUT.n722 0.0174092
R10227 VOUT.n716 VOUT.n713 0.0174092
R10228 VOUT.n707 VOUT.n704 0.0174092
R10229 VOUT.n698 VOUT.n695 0.0174092
R10230 VOUT.n689 VOUT.n686 0.0174092
R10231 VOUT.n680 VOUT.n677 0.0174092
R10232 VOUT.n671 VOUT.n668 0.0174092
R10233 VOUT.n662 VOUT.n659 0.0174092
R10234 VOUT.n653 VOUT.n650 0.0174092
R10235 VOUT.n644 VOUT.n641 0.0174092
R10236 VOUT.n635 VOUT.n632 0.0174092
R10237 VOUT.n626 VOUT.n623 0.0174092
R10238 VOUT.n617 VOUT.n614 0.0174092
R10239 VOUT.n608 VOUT.n605 0.0174092
R10240 VOUT.n599 VOUT.n596 0.0174092
R10241 VOUT.n590 VOUT.n587 0.0174092
R10242 VOUT.n581 VOUT.n578 0.0174092
R10243 VOUT.n572 VOUT.n569 0.0174092
R10244 VOUT.n940 VOUT.n937 0.0174092
R10245 VOUT.n931 VOUT.n928 0.0174092
R10246 VOUT.n922 VOUT.n919 0.0174092
R10247 VOUT.n913 VOUT.n910 0.0174092
R10248 VOUT.n904 VOUT.n901 0.0174092
R10249 VOUT.n895 VOUT.n892 0.0174092
R10250 VOUT.n886 VOUT.n883 0.0174092
R10251 VOUT.n877 VOUT.n874 0.0174092
R10252 VOUT.n868 VOUT.n865 0.0174092
R10253 VOUT.n859 VOUT.n856 0.0174092
R10254 VOUT.n850 VOUT.n847 0.0174092
R10255 VOUT.n841 VOUT.n838 0.0174092
R10256 VOUT.n832 VOUT.n829 0.0174092
R10257 VOUT.n823 VOUT.n820 0.0174092
R10258 VOUT.n814 VOUT.n811 0.0174092
R10259 VOUT.n805 VOUT.n802 0.0174092
R10260 VOUT.n796 VOUT.n793 0.0174092
R10261 VOUT.n787 VOUT.n784 0.0174092
R10262 VOUT.n778 VOUT.n775 0.0174092
R10263 VOUT.n769 VOUT.n766 0.0174092
R10264 VOUT.n760 VOUT.n757 0.0174092
R10265 VOUT.n1128 VOUT.n1125 0.0174092
R10266 VOUT.n1119 VOUT.n1116 0.0174092
R10267 VOUT.n1110 VOUT.n1107 0.0174092
R10268 VOUT.n1101 VOUT.n1098 0.0174092
R10269 VOUT.n1092 VOUT.n1089 0.0174092
R10270 VOUT.n1083 VOUT.n1080 0.0174092
R10271 VOUT.n1074 VOUT.n1071 0.0174092
R10272 VOUT.n1065 VOUT.n1062 0.0174092
R10273 VOUT.n1056 VOUT.n1053 0.0174092
R10274 VOUT.n1047 VOUT.n1044 0.0174092
R10275 VOUT.n1038 VOUT.n1035 0.0174092
R10276 VOUT.n1029 VOUT.n1026 0.0174092
R10277 VOUT.n1020 VOUT.n1017 0.0174092
R10278 VOUT.n1011 VOUT.n1008 0.0174092
R10279 VOUT.n1002 VOUT.n999 0.0174092
R10280 VOUT.n993 VOUT.n990 0.0174092
R10281 VOUT.n984 VOUT.n981 0.0174092
R10282 VOUT.n975 VOUT.n972 0.0174092
R10283 VOUT.n966 VOUT.n963 0.0174092
R10284 VOUT.n957 VOUT.n954 0.0174092
R10285 VOUT.n948 VOUT.n945 0.0174092
R10286 VOUT.n1316 VOUT.n1313 0.0174092
R10287 VOUT.n1307 VOUT.n1304 0.0174092
R10288 VOUT.n1298 VOUT.n1295 0.0174092
R10289 VOUT.n1289 VOUT.n1286 0.0174092
R10290 VOUT.n1280 VOUT.n1277 0.0174092
R10291 VOUT.n1271 VOUT.n1268 0.0174092
R10292 VOUT.n1262 VOUT.n1259 0.0174092
R10293 VOUT.n1253 VOUT.n1250 0.0174092
R10294 VOUT.n1244 VOUT.n1241 0.0174092
R10295 VOUT.n1235 VOUT.n1232 0.0174092
R10296 VOUT.n1226 VOUT.n1223 0.0174092
R10297 VOUT.n1217 VOUT.n1214 0.0174092
R10298 VOUT.n1208 VOUT.n1205 0.0174092
R10299 VOUT.n1199 VOUT.n1196 0.0174092
R10300 VOUT.n1190 VOUT.n1187 0.0174092
R10301 VOUT.n1181 VOUT.n1178 0.0174092
R10302 VOUT.n1172 VOUT.n1169 0.0174092
R10303 VOUT.n1163 VOUT.n1160 0.0174092
R10304 VOUT.n1154 VOUT.n1151 0.0174092
R10305 VOUT.n1145 VOUT.n1142 0.0174092
R10306 VOUT.n1136 VOUT.n1133 0.0174092
R10307 VOUT.n1504 VOUT.n1501 0.0174092
R10308 VOUT.n1495 VOUT.n1492 0.0174092
R10309 VOUT.n1486 VOUT.n1483 0.0174092
R10310 VOUT.n1477 VOUT.n1474 0.0174092
R10311 VOUT.n1468 VOUT.n1465 0.0174092
R10312 VOUT.n1459 VOUT.n1456 0.0174092
R10313 VOUT.n1450 VOUT.n1447 0.0174092
R10314 VOUT.n1441 VOUT.n1438 0.0174092
R10315 VOUT.n1432 VOUT.n1429 0.0174092
R10316 VOUT.n1423 VOUT.n1420 0.0174092
R10317 VOUT.n1414 VOUT.n1411 0.0174092
R10318 VOUT.n1405 VOUT.n1402 0.0174092
R10319 VOUT.n1396 VOUT.n1393 0.0174092
R10320 VOUT.n1387 VOUT.n1384 0.0174092
R10321 VOUT.n1378 VOUT.n1375 0.0174092
R10322 VOUT.n1369 VOUT.n1366 0.0174092
R10323 VOUT.n1360 VOUT.n1357 0.0174092
R10324 VOUT.n1351 VOUT.n1348 0.0174092
R10325 VOUT.n1342 VOUT.n1339 0.0174092
R10326 VOUT.n1333 VOUT.n1330 0.0174092
R10327 VOUT.n1324 VOUT.n1321 0.0174092
R10328 VOUT.n1692 VOUT.n1688 0.0174092
R10329 VOUT.n1683 VOUT.n1679 0.0174092
R10330 VOUT.n1674 VOUT.n1670 0.0174092
R10331 VOUT.n1665 VOUT.n1661 0.0174092
R10332 VOUT.n1656 VOUT.n1652 0.0174092
R10333 VOUT.n1647 VOUT.n1643 0.0174092
R10334 VOUT.n1638 VOUT.n1634 0.0174092
R10335 VOUT.n1629 VOUT.n1625 0.0174092
R10336 VOUT.n1620 VOUT.n1616 0.0174092
R10337 VOUT.n1611 VOUT.n1607 0.0174092
R10338 VOUT.n1602 VOUT.n1598 0.0174092
R10339 VOUT.n1593 VOUT.n1589 0.0174092
R10340 VOUT.n1584 VOUT.n1580 0.0174092
R10341 VOUT.n1575 VOUT.n1571 0.0174092
R10342 VOUT.n1566 VOUT.n1562 0.0174092
R10343 VOUT.n1557 VOUT.n1553 0.0174092
R10344 VOUT.n1548 VOUT.n1544 0.0174092
R10345 VOUT.n1539 VOUT.n1535 0.0174092
R10346 VOUT.n1530 VOUT.n1526 0.0174092
R10347 VOUT.n1521 VOUT.n1517 0.0174092
R10348 VOUT.n1512 VOUT.n1508 0.0174092
R10349 VOUT.n1880 VOUT.n1877 0.0174092
R10350 VOUT.n1871 VOUT.n1868 0.0174092
R10351 VOUT.n1862 VOUT.n1859 0.0174092
R10352 VOUT.n1853 VOUT.n1850 0.0174092
R10353 VOUT.n1844 VOUT.n1841 0.0174092
R10354 VOUT.n1835 VOUT.n1832 0.0174092
R10355 VOUT.n1826 VOUT.n1823 0.0174092
R10356 VOUT.n1817 VOUT.n1814 0.0174092
R10357 VOUT.n1808 VOUT.n1805 0.0174092
R10358 VOUT.n1799 VOUT.n1796 0.0174092
R10359 VOUT.n1790 VOUT.n1787 0.0174092
R10360 VOUT.n1781 VOUT.n1778 0.0174092
R10361 VOUT.n1772 VOUT.n1769 0.0174092
R10362 VOUT.n1763 VOUT.n1760 0.0174092
R10363 VOUT.n1754 VOUT.n1751 0.0174092
R10364 VOUT.n1745 VOUT.n1742 0.0174092
R10365 VOUT.n1736 VOUT.n1733 0.0174092
R10366 VOUT.n1727 VOUT.n1724 0.0174092
R10367 VOUT.n1718 VOUT.n1715 0.0174092
R10368 VOUT.n1709 VOUT.n1706 0.0174092
R10369 VOUT.n1700 VOUT.n1697 0.0174092
R10370 VOUT.n2068 VOUT.n2065 0.0174092
R10371 VOUT.n2059 VOUT.n2056 0.0174092
R10372 VOUT.n2050 VOUT.n2047 0.0174092
R10373 VOUT.n2041 VOUT.n2038 0.0174092
R10374 VOUT.n2032 VOUT.n2029 0.0174092
R10375 VOUT.n2023 VOUT.n2020 0.0174092
R10376 VOUT.n2014 VOUT.n2011 0.0174092
R10377 VOUT.n2005 VOUT.n2002 0.0174092
R10378 VOUT.n1996 VOUT.n1993 0.0174092
R10379 VOUT.n1987 VOUT.n1984 0.0174092
R10380 VOUT.n1978 VOUT.n1975 0.0174092
R10381 VOUT.n1969 VOUT.n1966 0.0174092
R10382 VOUT.n1960 VOUT.n1957 0.0174092
R10383 VOUT.n1951 VOUT.n1948 0.0174092
R10384 VOUT.n1942 VOUT.n1939 0.0174092
R10385 VOUT.n1933 VOUT.n1930 0.0174092
R10386 VOUT.n1924 VOUT.n1921 0.0174092
R10387 VOUT.n1915 VOUT.n1912 0.0174092
R10388 VOUT.n1906 VOUT.n1903 0.0174092
R10389 VOUT.n1897 VOUT.n1894 0.0174092
R10390 VOUT.n1888 VOUT.n1885 0.0174092
R10391 VOUT.n2256 VOUT.n2253 0.0174092
R10392 VOUT.n2247 VOUT.n2244 0.0174092
R10393 VOUT.n2238 VOUT.n2235 0.0174092
R10394 VOUT.n2229 VOUT.n2226 0.0174092
R10395 VOUT.n2220 VOUT.n2217 0.0174092
R10396 VOUT.n2211 VOUT.n2208 0.0174092
R10397 VOUT.n2202 VOUT.n2199 0.0174092
R10398 VOUT.n2193 VOUT.n2190 0.0174092
R10399 VOUT.n2184 VOUT.n2181 0.0174092
R10400 VOUT.n2175 VOUT.n2172 0.0174092
R10401 VOUT.n2166 VOUT.n2163 0.0174092
R10402 VOUT.n2157 VOUT.n2154 0.0174092
R10403 VOUT.n2148 VOUT.n2145 0.0174092
R10404 VOUT.n2139 VOUT.n2136 0.0174092
R10405 VOUT.n2130 VOUT.n2127 0.0174092
R10406 VOUT.n2121 VOUT.n2118 0.0174092
R10407 VOUT.n2112 VOUT.n2109 0.0174092
R10408 VOUT.n2103 VOUT.n2100 0.0174092
R10409 VOUT.n2094 VOUT.n2091 0.0174092
R10410 VOUT.n2085 VOUT.n2082 0.0174092
R10411 VOUT.n2076 VOUT.n2073 0.0174092
R10412 VOUT.n2264 VOUT.n2261 0.0174092
R10413 VOUT.n2271 VOUT.n2268 0.0174092
R10414 VOUT.n2278 VOUT.n2275 0.0174092
R10415 VOUT.n2285 VOUT.n2282 0.0174092
R10416 VOUT.n2292 VOUT.n2289 0.0174092
R10417 VOUT.n2299 VOUT.n2296 0.0174092
R10418 VOUT.n2306 VOUT.n2303 0.0174092
R10419 VOUT.n2313 VOUT.n2310 0.0174092
R10420 VOUT.n2320 VOUT.n2317 0.0174092
R10421 VOUT.n2327 VOUT.n2324 0.0174092
R10422 VOUT.n2334 VOUT.n2331 0.0174092
R10423 VOUT.n2341 VOUT.n2338 0.0174092
R10424 VOUT.n2348 VOUT.n2345 0.0174092
R10425 VOUT.n2355 VOUT.n2352 0.0174092
R10426 VOUT.n2362 VOUT.n2359 0.0174092
R10427 VOUT.n2369 VOUT.n2366 0.0174092
R10428 VOUT.n2376 VOUT.n2373 0.0174092
R10429 VOUT.n2383 VOUT.n2380 0.0174092
R10430 VOUT.n2390 VOUT.n2387 0.0174092
R10431 VOUT.n2397 VOUT.n2394 0.0174092
R10432 VOUT.n2404 VOUT.n2401 0.0174092
R10433 VOUT.n561 VOUT.n558 0.00635938
R10434 VOUT.n552 VOUT.n549 0.00635938
R10435 VOUT.n543 VOUT.n540 0.00635938
R10436 VOUT.n534 VOUT.n531 0.00635938
R10437 VOUT.n525 VOUT.n522 0.00635938
R10438 VOUT.n516 VOUT.n513 0.00635938
R10439 VOUT.n507 VOUT.n504 0.00635938
R10440 VOUT.n498 VOUT.n495 0.00635938
R10441 VOUT.n489 VOUT.n486 0.00635938
R10442 VOUT.n480 VOUT.n477 0.00635938
R10443 VOUT.n471 VOUT.n468 0.00635938
R10444 VOUT.n462 VOUT.n459 0.00635938
R10445 VOUT.n453 VOUT.n450 0.00635938
R10446 VOUT.n444 VOUT.n441 0.00635938
R10447 VOUT.n435 VOUT.n432 0.00635938
R10448 VOUT.n426 VOUT.n423 0.00635938
R10449 VOUT.n417 VOUT.n414 0.00635938
R10450 VOUT.n408 VOUT.n405 0.00635938
R10451 VOUT.n399 VOUT.n396 0.00635938
R10452 VOUT.n390 VOUT.n387 0.00635938
R10453 VOUT.n382 VOUT.n379 0.00635938
R10454 VOUT.n373 VOUT.n370 0.00635938
R10455 VOUT.n364 VOUT.n361 0.00635938
R10456 VOUT.n355 VOUT.n352 0.00635938
R10457 VOUT.n346 VOUT.n343 0.00635938
R10458 VOUT.n337 VOUT.n334 0.00635938
R10459 VOUT.n328 VOUT.n325 0.00635938
R10460 VOUT.n319 VOUT.n316 0.00635938
R10461 VOUT.n310 VOUT.n307 0.00635938
R10462 VOUT.n301 VOUT.n298 0.00635938
R10463 VOUT.n292 VOUT.n289 0.00635938
R10464 VOUT.n283 VOUT.n280 0.00635938
R10465 VOUT.n274 VOUT.n271 0.00635938
R10466 VOUT.n265 VOUT.n262 0.00635938
R10467 VOUT.n256 VOUT.n253 0.00635938
R10468 VOUT.n247 VOUT.n244 0.00635938
R10469 VOUT.n238 VOUT.n235 0.00635938
R10470 VOUT.n229 VOUT.n226 0.00635938
R10471 VOUT.n220 VOUT.n217 0.00635938
R10472 VOUT.n211 VOUT.n208 0.00635938
R10473 VOUT.n202 VOUT.n199 0.00635938
R10474 VOUT.n194 VOUT.n191 0.00635938
R10475 VOUT.n185 VOUT.n182 0.00635938
R10476 VOUT.n176 VOUT.n173 0.00635938
R10477 VOUT.n167 VOUT.n164 0.00635938
R10478 VOUT.n158 VOUT.n155 0.00635938
R10479 VOUT.n149 VOUT.n146 0.00635938
R10480 VOUT.n140 VOUT.n137 0.00635938
R10481 VOUT.n131 VOUT.n128 0.00635938
R10482 VOUT.n122 VOUT.n119 0.00635938
R10483 VOUT.n113 VOUT.n110 0.00635938
R10484 VOUT.n104 VOUT.n101 0.00635938
R10485 VOUT.n95 VOUT.n92 0.00635938
R10486 VOUT.n86 VOUT.n83 0.00635938
R10487 VOUT.n77 VOUT.n74 0.00635938
R10488 VOUT.n68 VOUT.n65 0.00635938
R10489 VOUT.n59 VOUT.n56 0.00635938
R10490 VOUT.n50 VOUT.n47 0.00635938
R10491 VOUT.n41 VOUT.n38 0.00635938
R10492 VOUT.n32 VOUT.n29 0.00635938
R10493 VOUT.n23 VOUT.n20 0.00635938
R10494 VOUT.n14 VOUT.n11 0.00635938
R10495 VOUT.n6 VOUT.n3 0.00635938
R10496 ndrv.n20 ndrv.t75 88.3811
R10497 ndrv.n2 ndrv.t67 88.1243
R10498 ndrv.n2 ndrv.t23 88.1243
R10499 ndrv.n2 ndrv.t119 88.1243
R10500 ndrv.n1 ndrv.t72 88.1243
R10501 ndrv.n1 ndrv.t30 88.1243
R10502 ndrv.n1 ndrv.t19 88.1243
R10503 ndrv.n1 ndrv.t101 88.1243
R10504 ndrv.n3 ndrv.t56 88.1243
R10505 ndrv.n3 ndrv.t28 88.1243
R10506 ndrv.n3 ndrv.t109 88.1243
R10507 ndrv.n3 ndrv.t97 88.1243
R10508 ndrv.n4 ndrv.t54 88.1243
R10509 ndrv.n4 ndrv.t50 88.1243
R10510 ndrv.n4 ndrv.t84 88.1243
R10511 ndrv.n4 ndrv.t49 88.1243
R10512 ndrv.n5 ndrv.t39 88.1243
R10513 ndrv.n5 ndrv.t117 88.1243
R10514 ndrv.n5 ndrv.t112 88.1243
R10515 ndrv.n5 ndrv.t27 88.1243
R10516 ndrv.n6 ndrv.t14 88.1243
R10517 ndrv.n6 ndrv.t5 88.1243
R10518 ndrv.n6 ndrv.t44 88.1243
R10519 ndrv.n6 ndrv.t51 88.1243
R10520 ndrv.n7 ndrv.t1 88.1243
R10521 ndrv.n7 ndrv.t6 88.1243
R10522 ndrv.n7 ndrv.t59 88.1243
R10523 ndrv.n7 ndrv.t110 88.1243
R10524 ndrv.n8 ndrv.t82 88.1243
R10525 ndrv.n8 ndrv.t48 88.1243
R10526 ndrv.n8 ndrv.t53 88.1243
R10527 ndrv.n8 ndrv.t95 88.1243
R10528 ndrv.n9 ndrv.t108 88.1243
R10529 ndrv.n9 ndrv.t25 88.1243
R10530 ndrv.n9 ndrv.t89 88.1243
R10531 ndrv.n9 ndrv.t98 88.1243
R10532 ndrv.n21 ndrv.t16 88.1243
R10533 ndrv.n21 ndrv.t12 88.1243
R10534 ndrv.n11 ndrv.t88 88.1243
R10535 ndrv.n11 ndrv.t58 88.1243
R10536 ndrv.n11 ndrv.t4 88.1243
R10537 ndrv.n11 ndrv.t0 88.1243
R10538 ndrv.n10 ndrv.t69 88.1243
R10539 ndrv.n10 ndrv.t47 88.1243
R10540 ndrv.n10 ndrv.t3 88.1243
R10541 ndrv.n10 ndrv.t76 88.1243
R10542 ndrv.n12 ndrv.t68 88.1243
R10543 ndrv.n12 ndrv.t24 88.1243
R10544 ndrv.n12 ndrv.t106 88.1243
R10545 ndrv.n12 ndrv.t73 88.1243
R10546 ndrv.n13 ndrv.t32 88.1243
R10547 ndrv.n13 ndrv.t21 88.1243
R10548 ndrv.n13 ndrv.t103 88.1243
R10549 ndrv.n13 ndrv.t92 88.1243
R10550 ndrv.n14 ndrv.t11 88.1243
R10551 ndrv.n14 ndrv.t91 88.1243
R10552 ndrv.n14 ndrv.t83 88.1243
R10553 ndrv.n14 ndrv.t43 88.1243
R10554 ndrv.n15 ndrv.t37 88.1243
R10555 ndrv.n15 ndrv.t71 88.1243
R10556 ndrv.n15 ndrv.t66 88.1243
R10557 ndrv.n15 ndrv.t60 88.1243
R10558 ndrv.n16 ndrv.t87 88.1243
R10559 ndrv.n16 ndrv.t96 88.1243
R10560 ndrv.n16 ndrv.t57 88.1243
R10561 ndrv.n16 ndrv.t61 88.1243
R10562 ndrv.n17 ndrv.t113 88.1243
R10563 ndrv.n17 ndrv.t33 88.1243
R10564 ndrv.n17 ndrv.t9 88.1243
R10565 ndrv.n17 ndrv.t90 88.1243
R10566 ndrv.n18 ndrv.t100 88.1243
R10567 ndrv.n18 ndrv.t18 88.1243
R10568 ndrv.n18 ndrv.t29 88.1243
R10569 ndrv.n18 ndrv.t70 88.1243
R10570 ndrv.n19 ndrv.t13 88.1243
R10571 ndrv.n19 ndrv.t22 88.1243
R10572 ndrv.n23 ndrv.t31 88.1243
R10573 ndrv.n23 ndrv.t20 88.1243
R10574 ndrv.n22 ndrv.t102 88.1243
R10575 ndrv.n22 ndrv.t63 88.1243
R10576 ndrv.n2 ndrv.t10 88.1243
R10577 ndrv.n2 ndrv.t7 88.1243
R10578 ndrv.n2 ndrv.t78 88.1243
R10579 ndrv.n2 ndrv.t55 88.1243
R10580 ndrv.n1 ndrv.t8 88.1243
R10581 ndrv.n1 ndrv.t85 88.1243
R10582 ndrv.n1 ndrv.t77 88.1243
R10583 ndrv.n1 ndrv.t38 88.1243
R10584 ndrv.n3 ndrv.t116 88.1243
R10585 ndrv.n3 ndrv.t81 88.1243
R10586 ndrv.n3 ndrv.t41 88.1243
R10587 ndrv.n3 ndrv.t35 88.1243
R10588 ndrv.n4 ndrv.t115 88.1243
R10589 ndrv.n4 ndrv.t107 88.1243
R10590 ndrv.n4 ndrv.t17 88.1243
R10591 ndrv.n4 ndrv.t105 88.1243
R10592 ndrv.n5 ndrv.t93 88.1243
R10593 ndrv.n5 ndrv.t52 88.1243
R10594 ndrv.n5 ndrv.t45 88.1243
R10595 ndrv.n5 ndrv.t80 88.1243
R10596 ndrv.n6 ndrv.t74 88.1243
R10597 ndrv.n6 ndrv.t64 88.1243
R10598 ndrv.n6 ndrv.t99 88.1243
R10599 ndrv.n6 ndrv.t111 88.1243
R10600 ndrv.n7 ndrv.t62 88.1243
R10601 ndrv.n7 ndrv.t65 88.1243
R10602 ndrv.n7 ndrv.t118 88.1243
R10603 ndrv.n7 ndrv.t42 88.1243
R10604 ndrv.n8 ndrv.t15 88.1243
R10605 ndrv.n8 ndrv.t104 88.1243
R10606 ndrv.n8 ndrv.t114 88.1243
R10607 ndrv.n8 ndrv.t34 88.1243
R10608 ndrv.n9 ndrv.t40 88.1243
R10609 ndrv.n9 ndrv.t79 88.1243
R10610 ndrv.n9 ndrv.t26 88.1243
R10611 ndrv.n9 ndrv.t36 88.1243
R10612 ndrv.n20 ndrv.t2 88.1243
R10613 ndrv.n20 ndrv.t46 88.1243
R10614 ndrv.n0 ndrv.t86 88.1243
R10615 ndrv.n0 ndrv.t94 88.1243
R10616 ndrv ndrv.n0 2.71641
R10617 ndrv.n9 ndrv.n24 3.26856
R10618 ndrv.n0 ndrv.n23 0.949823
R10619 ndrv.n23 ndrv.n21 0.807265
R10620 ndrv.n0 ndrv.n20 0.771066
R10621 ndrv.n17 ndrv.n18 0.687457
R10622 ndrv.n16 ndrv.n17 0.687457
R10623 ndrv.n15 ndrv.n16 0.687457
R10624 ndrv.n14 ndrv.n15 0.687457
R10625 ndrv.n13 ndrv.n14 0.687457
R10626 ndrv.n12 ndrv.n13 0.687457
R10627 ndrv.n10 ndrv.n12 0.687457
R10628 ndrv.n11 ndrv.n10 0.687457
R10629 ndrv.n21 ndrv.n11 0.687457
R10630 ndrv.n8 ndrv.n9 0.687457
R10631 ndrv.n7 ndrv.n8 0.687457
R10632 ndrv.n6 ndrv.n7 0.687457
R10633 ndrv.n5 ndrv.n6 0.687457
R10634 ndrv.n4 ndrv.n5 0.687457
R10635 ndrv.n3 ndrv.n4 0.687457
R10636 ndrv.n1 ndrv.n3 0.687457
R10637 ndrv.n2 ndrv.n1 0.687457
R10638 ndrv.n22 ndrv.n2 0.687457
R10639 ndrv.n23 ndrv.n22 0.579848
R10640 ndrv.n18 ndrv.n19 0.515717
R10641 VSS.n124 VSS.n123 292.505
R10642 VSS.n127 VSS.n126 292.5
R10643 VSS.n42 VSS.n41 292.5
R10644 VSS.n46 VSS.n45 292.5
R10645 VSS.n56 VSS.n55 292.5
R10646 VSS.n55 VSS.n54 292.5
R10647 VSS.n60 VSS.n59 292.5
R10648 VSS.n2873 VSS.n2872 292.5
R10649 VSS.n2866 VSS.n2865 292.5
R10650 VSS.n2859 VSS.n2858 292.5
R10651 VSS.n2852 VSS.n2851 292.5
R10652 VSS.n2845 VSS.n2844 292.5
R10653 VSS.n2835 VSS.n2834 292.5
R10654 VSS.n2828 VSS.n2827 292.5
R10655 VSS.n2821 VSS.n2820 292.5
R10656 VSS.n2819 VSS.n2818 292.5
R10657 VSS.n2812 VSS.n2811 292.5
R10658 VSS.n2805 VSS.n2804 292.5
R10659 VSS.n2798 VSS.n2797 292.5
R10660 VSS.n2791 VSS.n2790 292.5
R10661 VSS.n2784 VSS.n2783 292.5
R10662 VSS.n2777 VSS.n2776 292.5
R10663 VSS.n2770 VSS.n2769 292.5
R10664 VSS.n2764 VSS.n2763 292.5
R10665 VSS.n2756 VSS.n2755 292.5
R10666 VSS.n2749 VSS.n2748 292.5
R10667 VSS.n2742 VSS.n2741 292.5
R10668 VSS.n2735 VSS.n2734 292.5
R10669 VSS.n2728 VSS.n2727 292.5
R10670 VSS.n2721 VSS.n2720 292.5
R10671 VSS.n2711 VSS.n2710 292.5
R10672 VSS.n2704 VSS.n2703 292.5
R10673 VSS.n2697 VSS.n2696 292.5
R10674 VSS.n2695 VSS.n2694 292.5
R10675 VSS.n2688 VSS.n2687 292.5
R10676 VSS.n2681 VSS.n2680 292.5
R10677 VSS.n2674 VSS.n2673 292.5
R10678 VSS.n2667 VSS.n2666 292.5
R10679 VSS.n2660 VSS.n2659 292.5
R10680 VSS.n2653 VSS.n2652 292.5
R10681 VSS.n2646 VSS.n2645 292.5
R10682 VSS.n2640 VSS.n2639 292.5
R10683 VSS.n2632 VSS.n2631 292.5
R10684 VSS.n2625 VSS.n2624 292.5
R10685 VSS.n2618 VSS.n2617 292.5
R10686 VSS.n2611 VSS.n2610 292.5
R10687 VSS.n2604 VSS.n2603 292.5
R10688 VSS.n2597 VSS.n2596 292.5
R10689 VSS.n2587 VSS.n2586 292.5
R10690 VSS.n2580 VSS.n2579 292.5
R10691 VSS.n2573 VSS.n2572 292.5
R10692 VSS.n2571 VSS.n2570 292.5
R10693 VSS.n2564 VSS.n2563 292.5
R10694 VSS.n2557 VSS.n2556 292.5
R10695 VSS.n2550 VSS.n2549 292.5
R10696 VSS.n2543 VSS.n2542 292.5
R10697 VSS.n2536 VSS.n2535 292.5
R10698 VSS.n2529 VSS.n2528 292.5
R10699 VSS.n2522 VSS.n2521 292.5
R10700 VSS.n2516 VSS.n2515 292.5
R10701 VSS.n2508 VSS.n2507 292.5
R10702 VSS.n2501 VSS.n2500 292.5
R10703 VSS.n2494 VSS.n2493 292.5
R10704 VSS.n2487 VSS.n2486 292.5
R10705 VSS.n2480 VSS.n2479 292.5
R10706 VSS.n2473 VSS.n2472 292.5
R10707 VSS.n2463 VSS.n2462 292.5
R10708 VSS.n2456 VSS.n2455 292.5
R10709 VSS.n2449 VSS.n2448 292.5
R10710 VSS.n2446 VSS.n2445 292.5
R10711 VSS.n2440 VSS.n2439 292.5
R10712 VSS.n2433 VSS.n2432 292.5
R10713 VSS.n2426 VSS.n2425 292.5
R10714 VSS.n2419 VSS.n2418 292.5
R10715 VSS.n2412 VSS.n2411 292.5
R10716 VSS.n2405 VSS.n2404 292.5
R10717 VSS.n2398 VSS.n2397 292.5
R10718 VSS.n2392 VSS.n2391 292.5
R10719 VSS.n2384 VSS.n2383 292.5
R10720 VSS.n2377 VSS.n2376 292.5
R10721 VSS.n2370 VSS.n2369 292.5
R10722 VSS.n2363 VSS.n2362 292.5
R10723 VSS.n2356 VSS.n2355 292.5
R10724 VSS.n2349 VSS.n2348 292.5
R10725 VSS.n2339 VSS.n2338 292.5
R10726 VSS.n2332 VSS.n2331 292.5
R10727 VSS.n2325 VSS.n2324 292.5
R10728 VSS.n2322 VSS.n2321 292.5
R10729 VSS.n2316 VSS.n2315 292.5
R10730 VSS.n2309 VSS.n2308 292.5
R10731 VSS.n2302 VSS.n2301 292.5
R10732 VSS.n2295 VSS.n2294 292.5
R10733 VSS.n2288 VSS.n2287 292.5
R10734 VSS.n2281 VSS.n2280 292.5
R10735 VSS.n2877 VSS.n2876 292.5
R10736 VSS.n2245 VSS.n2244 292.5
R10737 VSS.n2278 VSS.n2277 292.5
R10738 VSS.n2284 VSS.n2283 292.5
R10739 VSS.n2290 VSS.n2289 292.5
R10740 VSS.n2298 VSS.n2297 292.5
R10741 VSS.n2304 VSS.n2303 292.5
R10742 VSS.n2312 VSS.n2311 292.5
R10743 VSS.n2318 VSS.n2317 292.5
R10744 VSS.n2328 VSS.n2327 292.5
R10745 VSS.n2334 VSS.n2333 292.5
R10746 VSS.n2342 VSS.n2341 292.5
R10747 VSS.n2347 VSS.n2346 292.5
R10748 VSS.n2353 VSS.n2352 292.5
R10749 VSS.n2361 VSS.n2360 292.5
R10750 VSS.n2367 VSS.n2366 292.5
R10751 VSS.n2375 VSS.n2374 292.5
R10752 VSS.n2381 VSS.n2380 292.5
R10753 VSS.n2389 VSS.n2388 292.5
R10754 VSS.n2396 VSS.n2395 292.5
R10755 VSS.n2402 VSS.n2401 292.5
R10756 VSS.n2408 VSS.n2407 292.5
R10757 VSS.n2414 VSS.n2413 292.5
R10758 VSS.n2422 VSS.n2421 292.5
R10759 VSS.n2428 VSS.n2427 292.5
R10760 VSS.n2436 VSS.n2435 292.5
R10761 VSS.n2442 VSS.n2441 292.5
R10762 VSS.n2452 VSS.n2451 292.5
R10763 VSS.n2458 VSS.n2457 292.5
R10764 VSS.n2466 VSS.n2465 292.5
R10765 VSS.n2471 VSS.n2470 292.5
R10766 VSS.n2477 VSS.n2476 292.5
R10767 VSS.n2485 VSS.n2484 292.5
R10768 VSS.n2491 VSS.n2490 292.5
R10769 VSS.n2499 VSS.n2498 292.5
R10770 VSS.n2505 VSS.n2504 292.5
R10771 VSS.n2513 VSS.n2512 292.5
R10772 VSS.n2520 VSS.n2519 292.5
R10773 VSS.n2526 VSS.n2525 292.5
R10774 VSS.n2532 VSS.n2531 292.5
R10775 VSS.n2538 VSS.n2537 292.5
R10776 VSS.n2546 VSS.n2545 292.5
R10777 VSS.n2552 VSS.n2551 292.5
R10778 VSS.n2560 VSS.n2559 292.5
R10779 VSS.n2566 VSS.n2565 292.5
R10780 VSS.n2576 VSS.n2575 292.5
R10781 VSS.n2582 VSS.n2581 292.5
R10782 VSS.n2590 VSS.n2589 292.5
R10783 VSS.n2595 VSS.n2594 292.5
R10784 VSS.n2601 VSS.n2600 292.5
R10785 VSS.n2609 VSS.n2608 292.5
R10786 VSS.n2615 VSS.n2614 292.5
R10787 VSS.n2623 VSS.n2622 292.5
R10788 VSS.n2629 VSS.n2628 292.5
R10789 VSS.n2637 VSS.n2636 292.5
R10790 VSS.n2644 VSS.n2643 292.5
R10791 VSS.n2650 VSS.n2649 292.5
R10792 VSS.n2656 VSS.n2655 292.5
R10793 VSS.n2662 VSS.n2661 292.5
R10794 VSS.n2670 VSS.n2669 292.5
R10795 VSS.n2676 VSS.n2675 292.5
R10796 VSS.n2684 VSS.n2683 292.5
R10797 VSS.n2690 VSS.n2689 292.5
R10798 VSS.n2700 VSS.n2699 292.5
R10799 VSS.n2706 VSS.n2705 292.5
R10800 VSS.n2714 VSS.n2713 292.5
R10801 VSS.n2719 VSS.n2718 292.5
R10802 VSS.n2725 VSS.n2724 292.5
R10803 VSS.n2733 VSS.n2732 292.5
R10804 VSS.n2739 VSS.n2738 292.5
R10805 VSS.n2747 VSS.n2746 292.5
R10806 VSS.n2753 VSS.n2752 292.5
R10807 VSS.n2761 VSS.n2760 292.5
R10808 VSS.n2768 VSS.n2767 292.5
R10809 VSS.n2774 VSS.n2773 292.5
R10810 VSS.n2780 VSS.n2779 292.5
R10811 VSS.n2786 VSS.n2785 292.5
R10812 VSS.n2794 VSS.n2793 292.5
R10813 VSS.n2800 VSS.n2799 292.5
R10814 VSS.n2808 VSS.n2807 292.5
R10815 VSS.n2814 VSS.n2813 292.5
R10816 VSS.n2824 VSS.n2823 292.5
R10817 VSS.n2830 VSS.n2829 292.5
R10818 VSS.n2838 VSS.n2837 292.5
R10819 VSS.n2843 VSS.n2842 292.5
R10820 VSS.n2849 VSS.n2848 292.5
R10821 VSS.n2857 VSS.n2856 292.5
R10822 VSS.n2863 VSS.n2862 292.5
R10823 VSS.n2871 VSS.n2870 292.5
R10824 VSS.n784 VSS.n783 292.5
R10825 VSS.n550 VSS.n549 292.5
R10826 VSS.n557 VSS.n556 292.5
R10827 VSS.n570 VSS.n569 292.5
R10828 VSS.n583 VSS.n582 292.5
R10829 VSS.n694 VSS.n693 292.5
R10830 VSS.n711 VSS.n710 292.5
R10831 VSS.n724 VSS.n723 292.5
R10832 VSS.n737 VSS.n736 292.5
R10833 VSS.n747 VSS.n746 292.5
R10834 VSS.n753 VSS.n752 292.5
R10835 VSS.n770 VSS.n769 292.5
R10836 VSS.n547 VSS.n546 292.5
R10837 VSS.n559 VSS.n558 292.5
R10838 VSS.n573 VSS.n572 292.5
R10839 VSS.n591 VSS.n590 292.5
R10840 VSS.n703 VSS.n702 292.5
R10841 VSS.n715 VSS.n714 292.5
R10842 VSS.n729 VSS.n728 292.5
R10843 VSS.n739 VSS.n738 292.5
R10844 VSS.n750 VSS.n749 292.5
R10845 VSS.n760 VSS.n759 292.5
R10846 VSS.n773 VSS.n772 292.5
R10847 VSS.n810 VSS.n809 292.5
R10848 VSS.n822 VSS.n821 292.5
R10849 VSS.n820 VSS.n819 292.5
R10850 VSS.n818 VSS.n817 292.5
R10851 VSS.n814 VSS.n813 292.5
R10852 VSS.n812 VSS.n811 292.5
R10853 VSS.n520 VSS.n519 292.5
R10854 VSS.n517 VSS.n516 292.5
R10855 VSS.n515 VSS.n514 292.5
R10856 VSS.n512 VSS.n511 292.5
R10857 VSS.n509 VSS.n508 292.5
R10858 VSS.n507 VSS.n506 292.5
R10859 VSS.n792 VSS.n791 292.5
R10860 VSS.n794 VSS.n793 292.5
R10861 VSS.n797 VSS.n796 292.5
R10862 VSS.n799 VSS.n798 292.5
R10863 VSS.n802 VSS.n801 292.5
R10864 VSS.n535 VSS.n534 292.5
R10865 VSS.n533 VSS.n532 292.5
R10866 VSS.n531 VSS.n530 292.5
R10867 VSS.n527 VSS.n526 292.5
R10868 VSS.n525 VSS.n524 292.5
R10869 VSS.n523 VSS.n522 292.5
R10870 VSS.n295 VSS.n294 292.5
R10871 VSS.n269 VSS.n268 292.5
R10872 VSS.n256 VSS.n255 292.5
R10873 VSS.n245 VSS.n244 292.5
R10874 VSS.n233 VSS.n232 292.5
R10875 VSS.n236 VSS.n235 292.5
R10876 VSS.n224 VSS.n223 292.5
R10877 VSS.n412 VSS.n411 292.5
R10878 VSS.n432 VSS.n431 292.5
R10879 VSS.n475 VSS.n474 292.5
R10880 VSS.n489 VSS.n488 292.5
R10881 VSS.n500 VSS.n499 292.5
R10882 VSS.n538 VSS.n537 292.5
R10883 VSS.n282 VSS.n281 292.5
R10884 VSS.n273 VSS.n272 292.5
R10885 VSS.n260 VSS.n259 292.5
R10886 VSS.n249 VSS.n248 292.5
R10887 VSS.n410 VSS.n409 292.5
R10888 VSS.n429 VSS.n428 292.5
R10889 VSS.n473 VSS.n472 292.5
R10890 VSS.n486 VSS.n485 292.5
R10891 VSS.n213 VSS.n212 292.5
R10892 VSS.n215 VSS.n214 292.5
R10893 VSS.n217 VSS.n216 292.5
R10894 VSS.n219 VSS.n218 292.5
R10895 VSS.n221 VSS.n220 292.5
R10896 VSS.n211 VSS.n210 292.5
R10897 VSS.n300 VSS.n299 292.5
R10898 VSS.n302 VSS.n301 292.5
R10899 VSS.n305 VSS.n304 292.5
R10900 VSS.n308 VSS.n307 292.5
R10901 VSS.n320 VSS.n319 292.5
R10902 VSS.n317 VSS.n316 292.5
R10903 VSS.n315 VSS.n314 292.5
R10904 VSS.n312 VSS.n311 292.5
R10905 VSS.n328 VSS.n327 292.5
R10906 VSS.n326 VSS.n325 292.5
R10907 VSS.n324 VSS.n323 292.5
R10908 VSS.n322 VSS.n321 292.5
R10909 VSS.n330 VSS.n329 292.5
R10910 VSS.n373 VSS.n359 292.5
R10911 VSS.n332 VSS.n331 292.5
R10912 VSS.n356 VSS.n355 292.5
R10913 VSS.n354 VSS.n353 292.5
R10914 VSS.n352 VSS.n351 292.5
R10915 VSS.n350 VSS.n349 292.5
R10916 VSS.n348 VSS.n347 292.5
R10917 VSS.n346 VSS.n345 292.5
R10918 VSS.n344 VSS.n343 292.5
R10919 VSS.n342 VSS.n341 292.5
R10920 VSS.n340 VSS.n339 292.5
R10921 VSS.n2247 VSS.n2246 292.5
R10922 VSS.n2249 VSS.n2248 292.5
R10923 VSS.n2251 VSS.n2250 292.5
R10924 VSS.n2253 VSS.n2252 292.5
R10925 VSS.n2255 VSS.n2254 292.5
R10926 VSS.n2257 VSS.n2256 292.5
R10927 VSS.n2259 VSS.n2258 292.5
R10928 VSS.n2261 VSS.n2260 292.5
R10929 VSS.n2263 VSS.n2262 292.5
R10930 VSS.n358 VSS.n357 292.5
R10931 VSS.n2268 VSS.n2267 292.5
R10932 VSS.n2273 VSS.n2272 292.5
R10933 VSS.n2271 VSS.n2270 292.5
R10934 VSS.n2921 VSS.n2920 292.5
R10935 VSS.n2924 VSS.n2923 292.5
R10936 VSS.n2928 VSS.n2927 292.5
R10937 VSS.n2932 VSS.n2931 292.5
R10938 VSS.n2936 VSS.n2935 292.5
R10939 VSS.n2940 VSS.n2939 292.5
R10940 VSS.n2943 VSS.n2942 292.5
R10941 VSS.n2947 VSS.n2946 292.5
R10942 VSS.n2951 VSS.n2950 292.5
R10943 VSS.n2955 VSS.n2954 292.5
R10944 VSS.n2959 VSS.n2958 292.5
R10945 VSS.n2963 VSS.n2962 292.5
R10946 VSS.n2967 VSS.n2966 292.5
R10947 VSS.n2971 VSS.n2970 292.5
R10948 VSS.n2984 VSS.n2983 292.5
R10949 VSS.n2988 VSS.n2987 292.5
R10950 VSS.n2993 VSS.n2992 292.5
R10951 VSS.n2998 VSS.n2997 292.5
R10952 VSS.n3002 VSS.n3001 292.5
R10953 VSS.n3007 VSS.n3006 292.5
R10954 VSS.n3011 VSS.n3010 292.5
R10955 VSS.n3013 VSS.n3012 292.5
R10956 VSS.n3018 VSS.n3017 292.5
R10957 VSS.n3022 VSS.n3021 292.5
R10958 VSS.n3027 VSS.n3026 292.5
R10959 VSS.n3031 VSS.n3030 292.5
R10960 VSS.n3036 VSS.n3035 292.5
R10961 VSS.n3040 VSS.n3039 292.5
R10962 VSS.n3045 VSS.n3044 292.5
R10963 VSS.n3050 VSS.n3049 292.5
R10964 VSS.n3054 VSS.n3053 292.5
R10965 VSS.n3059 VSS.n3058 292.5
R10966 VSS.n3063 VSS.n3062 292.5
R10967 VSS.n3068 VSS.n3067 292.5
R10968 VSS.n3072 VSS.n3071 292.5
R10969 VSS.n3077 VSS.n3076 292.5
R10970 VSS.n3081 VSS.n3080 292.5
R10971 VSS.n3086 VSS.n3085 292.5
R10972 VSS.n3090 VSS.n3089 292.5
R10973 VSS.n3092 VSS.n3091 292.5
R10974 VSS.n3097 VSS.n3096 292.5
R10975 VSS.n3101 VSS.n3100 292.5
R10976 VSS.n3106 VSS.n3105 292.5
R10977 VSS.n3110 VSS.n3109 292.5
R10978 VSS.n3115 VSS.n3114 292.5
R10979 VSS.n3119 VSS.n3118 292.5
R10980 VSS.n3124 VSS.n3123 292.5
R10981 VSS.n3129 VSS.n3128 292.5
R10982 VSS.n3133 VSS.n3132 292.5
R10983 VSS.n3138 VSS.n3137 292.5
R10984 VSS.n3142 VSS.n3141 292.5
R10985 VSS.n3147 VSS.n3146 292.5
R10986 VSS.n3151 VSS.n3150 292.5
R10987 VSS.n3156 VSS.n3155 292.5
R10988 VSS.n3160 VSS.n3159 292.5
R10989 VSS.n3165 VSS.n3164 292.5
R10990 VSS.n3169 VSS.n3168 292.5
R10991 VSS.n3171 VSS.n3170 292.5
R10992 VSS.n3176 VSS.n3175 292.5
R10993 VSS.n3180 VSS.n3179 292.5
R10994 VSS.n3185 VSS.n3184 292.5
R10995 VSS.n3189 VSS.n3188 292.5
R10996 VSS.n3194 VSS.n3193 292.5
R10997 VSS.n3198 VSS.n3197 292.5
R10998 VSS.n3203 VSS.n3202 292.5
R10999 VSS.n3208 VSS.n3207 292.5
R11000 VSS.n3212 VSS.n3211 292.5
R11001 VSS.n3217 VSS.n3216 292.5
R11002 VSS.n3221 VSS.n3220 292.5
R11003 VSS.n3226 VSS.n3225 292.5
R11004 VSS.n3230 VSS.n3229 292.5
R11005 VSS.n3235 VSS.n3234 292.5
R11006 VSS.n3239 VSS.n3238 292.5
R11007 VSS.n3244 VSS.n3243 292.5
R11008 VSS.n3248 VSS.n3247 292.5
R11009 VSS.n3250 VSS.n3249 292.5
R11010 VSS.n3255 VSS.n3254 292.5
R11011 VSS.n3259 VSS.n3258 292.5
R11012 VSS.n3264 VSS.n3263 292.5
R11013 VSS.n3268 VSS.n3267 292.5
R11014 VSS.n3273 VSS.n3272 292.5
R11015 VSS.n3277 VSS.n3276 292.5
R11016 VSS.n3282 VSS.n3281 292.5
R11017 VSS.n3287 VSS.n3286 292.5
R11018 VSS.n3291 VSS.n3290 292.5
R11019 VSS.n3296 VSS.n3295 292.5
R11020 VSS.n3300 VSS.n3299 292.5
R11021 VSS.n3305 VSS.n3304 292.5
R11022 VSS.n3309 VSS.n3308 292.5
R11023 VSS.n3314 VSS.n3313 292.5
R11024 VSS.n3318 VSS.n3317 292.5
R11025 VSS.n3323 VSS.n3322 292.5
R11026 VSS.n3327 VSS.n3326 292.5
R11027 VSS.n3329 VSS.n3328 292.5
R11028 VSS.n3334 VSS.n3333 292.5
R11029 VSS.n3338 VSS.n3337 292.5
R11030 VSS.n3343 VSS.n3342 292.5
R11031 VSS.n3347 VSS.n3346 292.5
R11032 VSS.n3352 VSS.n3351 292.5
R11033 VSS.n3356 VSS.n3355 292.5
R11034 VSS.n3363 VSS.n3362 292.5
R11035 VSS.n2914 VSS.n2913 292.5
R11036 VSS.n3447 VSS.n3446 292.5
R11037 VSS.n3373 VSS.n3372 292.5
R11038 VSS.n3378 VSS.n3377 292.5
R11039 VSS.n3377 VSS.n3376 292.5
R11040 VSS.n3383 VSS.n3382 292.5
R11041 VSS.n3382 VSS.n3381 292.5
R11042 VSS.n3388 VSS.n3387 292.5
R11043 VSS.n3387 VSS.n3386 292.5
R11044 VSS.n3393 VSS.n3392 292.5
R11045 VSS.n3392 VSS.n3391 292.5
R11046 VSS.n3398 VSS.n3397 292.5
R11047 VSS.n3397 VSS.n3396 292.5
R11048 VSS.n3403 VSS.n3402 292.5
R11049 VSS.n3402 VSS.n3401 292.5
R11050 VSS.n3408 VSS.n3407 292.5
R11051 VSS.n3407 VSS.n3406 292.5
R11052 VSS.n3413 VSS.n3412 292.5
R11053 VSS.n3412 VSS.n3411 292.5
R11054 VSS.n3418 VSS.n3417 292.5
R11055 VSS.n3417 VSS.n3416 292.5
R11056 VSS.n3423 VSS.n3422 292.5
R11057 VSS.n3422 VSS.n3421 292.5
R11058 VSS.n3428 VSS.n3427 292.5
R11059 VSS.n3427 VSS.n3426 292.5
R11060 VSS.n3433 VSS.n3432 292.5
R11061 VSS.n3432 VSS.n3431 292.5
R11062 VSS.n3438 VSS.n3437 292.5
R11063 VSS.n3437 VSS.n3436 292.5
R11064 VSS.n3443 VSS.n3442 292.5
R11065 VSS.n3442 VSS.n3441 292.5
R11066 VSS.n2895 VSS.n2894 292.5
R11067 VSS.n2893 VSS.n2892 292.5
R11068 VSS.n2891 VSS.n2890 292.5
R11069 VSS.n2889 VSS.n2888 292.5
R11070 VSS.n2887 VSS.n2886 292.5
R11071 VSS.n2885 VSS.n2884 292.5
R11072 VSS.n2883 VSS.n2882 292.5
R11073 VSS.n2881 VSS.n2880 292.5
R11074 VSS.n129 VSS.n128 292.5
R11075 VSS.n131 VSS.n130 292.5
R11076 VSS.n133 VSS.n132 292.5
R11077 VSS.n135 VSS.n134 292.5
R11078 VSS.n137 VSS.n136 292.5
R11079 VSS.n139 VSS.n138 292.5
R11080 VSS.n141 VSS.n140 292.5
R11081 VSS.n143 VSS.n142 292.5
R11082 VSS.n145 VSS.n144 292.5
R11083 VSS.n147 VSS.n146 292.5
R11084 VSS.n2897 VSS.n2896 292.5
R11085 VSS.n110 VSS.n109 292.5
R11086 VSS.n115 VSS.n114 292.5
R11087 VSS.n64 VSS.n63 292.5
R11088 VSS.n85 VSS.n84 292.5
R11089 VSS.n90 VSS.n89 292.5
R11090 VSS.n104 VSS.n103 292.5
R11091 VSS.n100 VSS.n99 292.5
R11092 VSS.n96 VSS.n95 292.5
R11093 VSS.n94 VSS.n93 292.5
R11094 VSS.n112 VSS.n111 292.5
R11095 VSS.n117 VSS.n116 292.5
R11096 VSS.n120 VSS.n119 292.5
R11097 VSS.n122 VSS.n121 292.5
R11098 VSS.n152 VSS.n151 292.5
R11099 VSS.n76 VSS.n75 292.5
R11100 VSS.n73 VSS.n72 292.5
R11101 VSS.n62 VSS.n61 292.5
R11102 VSS.n58 VSS.n57 292.5
R11103 VSS.n53 VSS.n52 292.5
R11104 VSS.n52 VSS.n51 292.5
R11105 VSS.n49 VSS.n48 292.5
R11106 VSS.n1477 VSS.n1476 292.5
R11107 VSS.n1469 VSS.n1468 292.5
R11108 VSS.n1471 VSS.n1470 292.5
R11109 VSS.n1473 VSS.n1472 292.5
R11110 VSS.n1475 VSS.n1474 292.5
R11111 VSS.n1467 VSS.n1466 292.5
R11112 VSS.n1357 VSS.n1356 292.5
R11113 VSS.n1349 VSS.n1348 292.5
R11114 VSS.n1351 VSS.n1350 292.5
R11115 VSS.n1353 VSS.n1352 292.5
R11116 VSS.n1355 VSS.n1354 292.5
R11117 VSS.n1347 VSS.n1346 292.5
R11118 VSS.n1234 VSS.n1233 292.5
R11119 VSS.n1226 VSS.n1225 292.5
R11120 VSS.n1228 VSS.n1227 292.5
R11121 VSS.n1230 VSS.n1229 292.5
R11122 VSS.n1232 VSS.n1231 292.5
R11123 VSS.n1224 VSS.n1223 292.5
R11124 VSS.n1131 VSS.n1130 292.5
R11125 VSS.n1123 VSS.n1122 292.5
R11126 VSS.n1125 VSS.n1124 292.5
R11127 VSS.n1127 VSS.n1126 292.5
R11128 VSS.n1129 VSS.n1128 292.5
R11129 VSS.n1121 VSS.n1120 292.5
R11130 VSS.n1000 VSS.n999 292.5
R11131 VSS.n992 VSS.n991 292.5
R11132 VSS.n994 VSS.n993 292.5
R11133 VSS.n996 VSS.n995 292.5
R11134 VSS.n998 VSS.n997 292.5
R11135 VSS.n990 VSS.n989 292.5
R11136 VSS.n681 VSS.n680 292.5
R11137 VSS.n673 VSS.n672 292.5
R11138 VSS.n675 VSS.n674 292.5
R11139 VSS.n677 VSS.n676 292.5
R11140 VSS.n679 VSS.n678 292.5
R11141 VSS.n671 VSS.n670 292.5
R11142 VSS.n807 VSS.n806 292.5
R11143 VSS.n804 VSS.n803 292.5
R11144 VSS.n659 VSS.n658 292.5
R11145 VSS.n663 VSS.n662 292.5
R11146 VSS.n668 VSS.n667 292.5
R11147 VSS.n665 VSS.n664 292.5
R11148 VSS.n978 VSS.n977 292.5
R11149 VSS.n982 VSS.n981 292.5
R11150 VSS.n987 VSS.n986 292.5
R11151 VSS.n984 VSS.n983 292.5
R11152 VSS.n1109 VSS.n1108 292.5
R11153 VSS.n1112 VSS.n1111 292.5
R11154 VSS.n1118 VSS.n1117 292.5
R11155 VSS.n1114 VSS.n1113 292.5
R11156 VSS.n1212 VSS.n1211 292.5
R11157 VSS.n1216 VSS.n1215 292.5
R11158 VSS.n1221 VSS.n1220 292.5
R11159 VSS.n1218 VSS.n1217 292.5
R11160 VSS.n1338 VSS.n1337 292.5
R11161 VSS.n1341 VSS.n1340 292.5
R11162 VSS.n1344 VSS.n1343 292.5
R11163 VSS.n2 VSS.n1 292.5
R11164 VSS.n4 VSS.n3 292.5
R11165 VSS.n7 VSS.n6 292.5
R11166 VSS.n11 VSS.n10 292.5
R11167 VSS.n14 VSS.n13 292.5
R11168 VSS.n16 VSS.n15 292.5
R11169 VSS.n19 VSS.n18 292.5
R11170 VSS.n25 VSS.n24 292.5
R11171 VSS.n28 VSS.n27 292.5
R11172 VSS.n30 VSS.n29 292.5
R11173 VSS.n36 VSS.n35 292.5
R11174 VSS.n1584 VSS.n1583 292.5
R11175 VSS.n1586 VSS.n1585 292.5
R11176 VSS.n1588 VSS.n1587 292.5
R11177 VSS.n1590 VSS.n1589 292.5
R11178 VSS.n1592 VSS.n1591 292.5
R11179 VSS.n21 VSS.n20 292.5
R11180 VSS.n825 VSS.n824 292.5
R11181 VSS.n836 VSS.n835 292.5
R11182 VSS.n849 VSS.n848 292.5
R11183 VSS.n862 VSS.n861 292.5
R11184 VSS.n873 VSS.n872 292.5
R11185 VSS.n884 VSS.n883 292.5
R11186 VSS.n686 VSS.n685 292.5
R11187 VSS.n689 VSS.n688 292.5
R11188 VSS.n894 VSS.n893 292.5
R11189 VSS.n909 VSS.n908 292.5
R11190 VSS.n951 VSS.n950 292.5
R11191 VSS.n963 VSS.n962 292.5
R11192 VSS.n976 VSS.n975 292.5
R11193 VSS.n1010 VSS.n1009 292.5
R11194 VSS.n1012 VSS.n1011 292.5
R11195 VSS.n1030 VSS.n1029 292.5
R11196 VSS.n1044 VSS.n1043 292.5
R11197 VSS.n1055 VSS.n1054 292.5
R11198 VSS.n1098 VSS.n1097 292.5
R11199 VSS.n1134 VSS.n1133 292.5
R11200 VSS.n1145 VSS.n1144 292.5
R11201 VSS.n1152 VSS.n1151 292.5
R11202 VSS.n1164 VSS.n1163 292.5
R11203 VSS.n1175 VSS.n1174 292.5
R11204 VSS.n1187 VSS.n1186 292.5
R11205 VSS.n1201 VSS.n1200 292.5
R11206 VSS.n1239 VSS.n1238 292.5
R11207 VSS.n1281 VSS.n1280 292.5
R11208 VSS.n1294 VSS.n1293 292.5
R11209 VSS.n1306 VSS.n1305 292.5
R11210 VSS.n1316 VSS.n1315 292.5
R11211 VSS.n1323 VSS.n1322 292.5
R11212 VSS.n1360 VSS.n1359 292.5
R11213 VSS.n1370 VSS.n1369 292.5
R11214 VSS.n1382 VSS.n1381 292.5
R11215 VSS.n1424 VSS.n1423 292.5
R11216 VSS.n1437 VSS.n1436 292.5
R11217 VSS.n1456 VSS.n1455 292.5
R11218 VSS.n1459 VSS.n1458 292.5
R11219 VSS.n1481 VSS.n1480 292.5
R11220 VSS.n1491 VSS.n1490 292.5
R11221 VSS.n1504 VSS.n1503 292.5
R11222 VSS.n1514 VSS.n1513 292.5
R11223 VSS.n1530 VSS.n1529 292.5
R11224 VSS.n1575 VSS.n1574 292.5
R11225 VSS.n1596 VSS.n1595 292.5
R11226 VSS.n1605 VSS.n1604 292.5
R11227 VSS.n1617 VSS.n1616 292.5
R11228 VSS.n1619 VSS.n1618 292.5
R11229 VSS.n1641 VSS.n1640 292.5
R11230 VSS.n1655 VSS.n1654 292.5
R11231 VSS.n846 VSS.n845 292.5
R11232 VSS.n859 VSS.n858 292.5
R11233 VSS.n870 VSS.n869 292.5
R11234 VSS.n882 VSS.n881 292.5
R11235 VSS.n901 VSS.n900 292.5
R11236 VSS.n943 VSS.n942 292.5
R11237 VSS.n954 VSS.n953 292.5
R11238 VSS.n967 VSS.n966 292.5
R11239 VSS.n1021 VSS.n1020 292.5
R11240 VSS.n1034 VSS.n1033 292.5
R11241 VSS.n1047 VSS.n1046 292.5
R11242 VSS.n1063 VSS.n1062 292.5
R11243 VSS.n1155 VSS.n1154 292.5
R11244 VSS.n1167 VSS.n1166 292.5
R11245 VSS.n1177 VSS.n1176 292.5
R11246 VSS.n1192 VSS.n1191 292.5
R11247 VSS.n1284 VSS.n1283 292.5
R11248 VSS.n1298 VSS.n1297 292.5
R11249 VSS.n1308 VSS.n1307 292.5
R11250 VSS.n1320 VSS.n1319 292.5
R11251 VSS.n1379 VSS.n1378 292.5
R11252 VSS.n1422 VSS.n1421 292.5
R11253 VSS.n1434 VSS.n1433 292.5
R11254 VSS.n1448 VSS.n1447 292.5
R11255 VSS.n1489 VSS.n1488 292.5
R11256 VSS.n1502 VSS.n1501 292.5
R11257 VSS.n1523 VSS.n1522 292.5
R11258 VSS.n1566 VSS.n1565 292.5
R11259 VSS.n1608 VSS.n1607 292.5
R11260 VSS.n1624 VSS.n1623 292.5
R11261 VSS.n1632 VSS.n1631 292.5
R11262 VSS.n1645 VSS.n1644 292.5
R11263 VSS.n881 VSS.n880 270.034
R11264 VSS.n248 VSS.n247 270.034
R11265 VSS.n311 VSS.n310 270.034
R11266 VSS.n1607 VSS.n1606 270.034
R11267 VSS.n24 VSS.n23 270.034
R11268 VSS.n10 VSS.n9 270.034
R11269 VSS.n1447 VSS.n1446 270.034
R11270 VSS.n1343 VSS.n1342 270.034
R11271 VSS.n1319 VSS.n1318 270.034
R11272 VSS.n1154 VSS.n1153 270.034
R11273 VSS.n1191 VSS.n1190 270.034
R11274 VSS.n1117 VSS.n1115 270.034
R11275 VSS.n1215 VSS.n1214 270.034
R11276 VSS.n1020 VSS.n1019 270.034
R11277 VSS.n981 VSS.n980 270.034
R11278 VSS.n662 VSS.n661 270.034
R11279 VSS.n372 VSS.n360 161.944
R11280 VSS.n335 VSS.n334 161.944
R11281 VSS.n372 VSS.n371 161.944
R11282 VSS.n2912 VSS.n2911 161.944
R11283 VSS.n2266 VSS.n2265 140.44
R11284 VSS.n530 VSS.n529 132.531
R11285 VSS.n817 VSS.n816 127.334
R11286 VSS.n41 VSS.n40 117.719
R11287 VSS.n114 VSS.n113 117.719
R11288 VSS.n3017 VSS.n3016 117.719
R11289 VSS.n3026 VSS.n3025 117.719
R11290 VSS.n3035 VSS.n3034 117.719
R11291 VSS.n3044 VSS.n3043 117.719
R11292 VSS.n3096 VSS.n3095 117.719
R11293 VSS.n3105 VSS.n3104 117.719
R11294 VSS.n3114 VSS.n3113 117.719
R11295 VSS.n3123 VSS.n3122 117.719
R11296 VSS.n3175 VSS.n3174 117.719
R11297 VSS.n3184 VSS.n3183 117.719
R11298 VSS.n3193 VSS.n3192 117.719
R11299 VSS.n3202 VSS.n3201 117.719
R11300 VSS.n3254 VSS.n3253 117.719
R11301 VSS.n3263 VSS.n3262 117.719
R11302 VSS.n3272 VSS.n3271 117.719
R11303 VSS.n3281 VSS.n3280 117.719
R11304 VSS.n3333 VSS.n3332 117.719
R11305 VSS.n3342 VSS.n3341 117.719
R11306 VSS.n3351 VSS.n3350 117.719
R11307 VSS.n3362 VSS.n3361 117.719
R11308 VSS.n2280 VSS.n2279 117.719
R11309 VSS.n2294 VSS.n2293 117.719
R11310 VSS.n2308 VSS.n2307 117.719
R11311 VSS.n2391 VSS.n2390 117.719
R11312 VSS.n2404 VSS.n2403 117.719
R11313 VSS.n2418 VSS.n2417 117.719
R11314 VSS.n2432 VSS.n2431 117.719
R11315 VSS.n2515 VSS.n2514 117.719
R11316 VSS.n2528 VSS.n2527 117.719
R11317 VSS.n2542 VSS.n2541 117.719
R11318 VSS.n2556 VSS.n2555 117.719
R11319 VSS.n2570 VSS.n2569 117.719
R11320 VSS.n2639 VSS.n2638 117.719
R11321 VSS.n2652 VSS.n2651 117.719
R11322 VSS.n2666 VSS.n2665 117.719
R11323 VSS.n2680 VSS.n2679 117.719
R11324 VSS.n2694 VSS.n2693 117.719
R11325 VSS.n2763 VSS.n2762 117.719
R11326 VSS.n2776 VSS.n2775 117.719
R11327 VSS.n2790 VSS.n2789 117.719
R11328 VSS.n2804 VSS.n2803 117.719
R11329 VSS.n2818 VSS.n2817 117.719
R11330 VSS.n2865 VSS.n2864 117.719
R11331 VSS.n2851 VSS.n2850 117.719
R11332 VSS.n2834 VSS.n2833 117.719
R11333 VSS.n2755 VSS.n2754 117.719
R11334 VSS.n2741 VSS.n2740 117.719
R11335 VSS.n2727 VSS.n2726 117.719
R11336 VSS.n2710 VSS.n2709 117.719
R11337 VSS.n2631 VSS.n2630 117.719
R11338 VSS.n2617 VSS.n2616 117.719
R11339 VSS.n2603 VSS.n2602 117.719
R11340 VSS.n2586 VSS.n2585 117.719
R11341 VSS.n2507 VSS.n2506 117.719
R11342 VSS.n2493 VSS.n2492 117.719
R11343 VSS.n2479 VSS.n2478 117.719
R11344 VSS.n2462 VSS.n2461 117.719
R11345 VSS.n2448 VSS.n2447 117.719
R11346 VSS.n2383 VSS.n2382 117.719
R11347 VSS.n2369 VSS.n2368 117.719
R11348 VSS.n2355 VSS.n2354 117.719
R11349 VSS.n2338 VSS.n2337 117.719
R11350 VSS.n2324 VSS.n2323 117.719
R11351 VSS.n2997 VSS.n2996 117.719
R11352 VSS.n3006 VSS.n3005 117.719
R11353 VSS.n3049 VSS.n3048 117.719
R11354 VSS.n3058 VSS.n3057 117.719
R11355 VSS.n3067 VSS.n3066 117.719
R11356 VSS.n3076 VSS.n3075 117.719
R11357 VSS.n3085 VSS.n3084 117.719
R11358 VSS.n3128 VSS.n3127 117.719
R11359 VSS.n3137 VSS.n3136 117.719
R11360 VSS.n3146 VSS.n3145 117.719
R11361 VSS.n3155 VSS.n3154 117.719
R11362 VSS.n3164 VSS.n3163 117.719
R11363 VSS.n3207 VSS.n3206 117.719
R11364 VSS.n3216 VSS.n3215 117.719
R11365 VSS.n3225 VSS.n3224 117.719
R11366 VSS.n3234 VSS.n3233 117.719
R11367 VSS.n3243 VSS.n3242 117.719
R11368 VSS.n3286 VSS.n3285 117.719
R11369 VSS.n3295 VSS.n3294 117.719
R11370 VSS.n3304 VSS.n3303 117.719
R11371 VSS.n3313 VSS.n3312 117.719
R11372 VSS.n3322 VSS.n3321 117.719
R11373 VSS.n373 VSS.n338 105.766
R11374 VSS.n373 VSS.n372 105.766
R11375 VSS.n373 VSS.n335 105.766
R11376 VSS.n2268 VSS.n2266 105.766
R11377 VSS.n2914 VSS.n2912 105.766
R11378 VSS.n32 VSS.n31 105.766
R11379 VSS.n371 VSS.n370 105.766
R11380 VSS.n2911 VSS.n2910 105.766
R11381 VSS.n78 VSS.n77 105.766
R11382 VSS.n34 VSS.n33 105.766
R11383 VSS.n1622 VSS.n1621 105.766
R11384 VSS.n2910 VSS.n2909 98.0106
R11385 VSS.n304 VSS.n303 93.9796
R11386 VSS.n2983 VSS.n2982 90.6381
R11387 VSS.n2992 VSS.n2991 90.6381
R11388 VSS.n40 VSS.n39 87.3927
R11389 VSS.n3361 VSS.n3360 87.3925
R11390 VSS.n2346 VSS.n2345 80.9725
R11391 VSS.n2360 VSS.n2359 80.9725
R11392 VSS.n2374 VSS.n2373 80.9725
R11393 VSS.n2388 VSS.n2387 80.9725
R11394 VSS.n2470 VSS.n2469 80.9725
R11395 VSS.n2484 VSS.n2483 80.9725
R11396 VSS.n2498 VSS.n2497 80.9725
R11397 VSS.n2512 VSS.n2511 80.9725
R11398 VSS.n2594 VSS.n2593 80.9725
R11399 VSS.n2608 VSS.n2607 80.9725
R11400 VSS.n2622 VSS.n2621 80.9725
R11401 VSS.n2636 VSS.n2635 80.9725
R11402 VSS.n2718 VSS.n2717 80.9725
R11403 VSS.n2732 VSS.n2731 80.9725
R11404 VSS.n2746 VSS.n2745 80.9725
R11405 VSS.n2760 VSS.n2759 80.9725
R11406 VSS.n2842 VSS.n2841 80.9725
R11407 VSS.n2856 VSS.n2855 80.9725
R11408 VSS.n2870 VSS.n2869 80.9725
R11409 VSS.n736 VSS.n735 80.9725
R11410 VSS.n268 VSS.n267 80.9725
R11411 VSS.n244 VSS.n243 80.9725
R11412 VSS.n235 VSS.n234 80.9725
R11413 VSS.n281 VSS.n280 80.9725
R11414 VSS.n319 VSS.n318 80.9725
R11415 VSS.n338 VSS.n336 80.9725
R11416 VSS.n2912 VSS.n2898 80.9725
R11417 VSS.n2837 VSS.n2836 80.9721
R11418 VSS.n2823 VSS.n2822 80.9721
R11419 VSS.n2807 VSS.n2806 80.9721
R11420 VSS.n2793 VSS.n2792 80.9721
R11421 VSS.n2779 VSS.n2778 80.9721
R11422 VSS.n2713 VSS.n2712 80.9721
R11423 VSS.n2699 VSS.n2698 80.9721
R11424 VSS.n2683 VSS.n2682 80.9721
R11425 VSS.n2669 VSS.n2668 80.9721
R11426 VSS.n2655 VSS.n2654 80.9721
R11427 VSS.n2589 VSS.n2588 80.9721
R11428 VSS.n2575 VSS.n2574 80.9721
R11429 VSS.n2559 VSS.n2558 80.9721
R11430 VSS.n2545 VSS.n2544 80.9721
R11431 VSS.n2531 VSS.n2530 80.9721
R11432 VSS.n2465 VSS.n2464 80.9721
R11433 VSS.n2451 VSS.n2450 80.9721
R11434 VSS.n2435 VSS.n2434 80.9721
R11435 VSS.n2421 VSS.n2420 80.9721
R11436 VSS.n2407 VSS.n2406 80.9721
R11437 VSS.n2341 VSS.n2340 80.9721
R11438 VSS.n2327 VSS.n2326 80.9721
R11439 VSS.n2311 VSS.n2310 80.9721
R11440 VSS.n2297 VSS.n2296 80.9721
R11441 VSS.n2283 VSS.n2282 80.9721
R11442 VSS.n723 VSS.n722 80.9721
R11443 VSS.n693 VSS.n692 80.9721
R11444 VSS.n569 VSS.n568 80.9721
R11445 VSS.n488 VSS.n487 80.9721
R11446 VSS.n431 VSS.n430 80.9721
R11447 VSS.n338 VSS.n337 80.9721
R11448 VSS.n2266 VSS.n2264 80.9721
R11449 VSS.n858 VSS.n857 80.9719
R11450 VSS.n848 VSS.n847 80.9719
R11451 VSS.n872 VSS.n871 80.9719
R11452 VSS.n685 VSS.n684 80.9719
R11453 VSS.n893 VSS.n892 80.9719
R11454 VSS.n975 VSS.n974 80.9719
R11455 VSS.n1043 VSS.n1042 80.9719
R11456 VSS.n1144 VSS.n1143 80.9719
R11457 VSS.n1163 VSS.n1162 80.9719
R11458 VSS.n1186 VSS.n1185 80.9719
R11459 VSS.n1238 VSS.n1237 80.9719
R11460 VSS.n1293 VSS.n1292 80.9719
R11461 VSS.n1381 VSS.n1380 80.9719
R11462 VSS.n1436 VSS.n1435 80.9719
R11463 VSS.n1458 VSS.n1457 80.9719
R11464 VSS.n1513 VSS.n1512 80.9719
R11465 VSS.n1604 VSS.n1603 80.9719
R11466 VSS.n1654 VSS.n1653 80.9719
R11467 VSS.n84 VSS.n83 80.9719
R11468 VSS.n103 VSS.n102 80.9719
R11469 VSS.n119 VSS.n118 80.9719
R11470 VSS.n151 VSS.n150 80.9719
R11471 VSS.n796 VSS.n795 80.9719
R11472 VSS.n801 VSS.n800 80.9719
R11473 VSS.n248 VSS.n246 80.9719
R11474 VSS.n428 VSS.n427 80.9719
R11475 VSS.n485 VSS.n484 80.9719
R11476 VSS.n702 VSS.n701 80.9719
R11477 VSS.n728 VSS.n727 80.9719
R11478 VSS.n749 VSS.n748 80.9719
R11479 VSS.n772 VSS.n771 80.9719
R11480 VSS.n511 VSS.n510 80.9719
R11481 VSS.n314 VSS.n313 80.9719
R11482 VSS.n99 VSS.n98 80.9719
R11483 VSS.n93 VSS.n92 80.9719
R11484 VSS.n1623 VSS.n1622 80.9719
R11485 VSS.n1644 VSS.n1643 80.9719
R11486 VSS.n77 VSS.n73 80.9719
R11487 VSS.n77 VSS.n76 80.9719
R11488 VSS.n27 VSS.n26 80.9719
R11489 VSS.n35 VSS.n34 80.9719
R11490 VSS.n13 VSS.n12 80.9719
R11491 VSS.n18 VSS.n17 80.9719
R11492 VSS.n1501 VSS.n1500 80.9719
R11493 VSS.n1447 VSS.n1445 80.9719
R11494 VSS.n1 VSS.n0 80.9719
R11495 VSS.n6 VSS.n5 80.9719
R11496 VSS.n1340 VSS.n1339 80.9719
R11497 VSS.n1297 VSS.n1296 80.9719
R11498 VSS.n1319 VSS.n1317 80.9719
R11499 VSS.n1166 VSS.n1165 80.9719
R11500 VSS.n1191 VSS.n1189 80.9719
R11501 VSS.n1215 VSS.n1213 80.9719
R11502 VSS.n1111 VSS.n1110 80.9719
R11503 VSS.n1033 VSS.n1032 80.9719
R11504 VSS.n1062 VSS.n1061 80.9719
R11505 VSS.n966 VSS.n965 80.9719
R11506 VSS.n981 VSS.n979 80.9719
R11507 VSS.n662 VSS.n660 80.9719
R11508 VSS.n806 VSS.n805 80.9719
R11509 VSS.n667 VSS.n666 80.9719
R11510 VSS.n986 VSS.n985 80.9719
R11511 VSS.n1117 VSS.n1116 80.9719
R11512 VSS.n1220 VSS.n1219 80.9719
R11513 VSS.n908 VSS.n907 80.9719
R11514 VSS.n1009 VSS.n1008 80.9719
R11515 VSS.n1054 VSS.n1053 80.9719
R11516 VSS.n1305 VSS.n1304 80.9719
R11517 VSS.n1322 VSS.n1321 80.9719
R11518 VSS.n1480 VSS.n1479 80.9719
R11519 VSS.n1529 VSS.n1528 80.9719
R11520 VSS.n1616 VSS.n1615 80.9719
R11521 VSS.n869 VSS.n868 80.9719
R11522 VSS.n900 VSS.n899 80.9719
R11523 VSS.n1378 VSS.n1377 80.9719
R11524 VSS.n1522 VSS.n1521 80.9719
R11525 VSS.n2909 VSS.n2908 75.1416
R11526 VSS.n3360 VSS.n3359 75.1416
R11527 VSS.n370 VSS.n369 64.6872
R11528 VSS.n2910 VSS.n2907 64.6872
R11529 VSS.n307 VSS.n306 59.4692
R11530 VSS.n2244 VSS.n2243 59.4689
R11531 VSS.n499 VSS.n498 59.4689
R11532 VSS.n549 VSS.n548 59.4689
R11533 VSS.n752 VSS.n751 59.4689
R11534 VSS.n783 VSS.n782 59.4689
R11535 VSS.n519 VSS.n518 59.4689
R11536 VSS.n514 VSS.n513 59.4689
R11537 VSS.n299 VSS.n298 59.4689
R11538 VSS.n546 VSS.n545 59.4689
R11539 VSS.n572 VSS.n571 59.4689
R11540 VSS.n322 VSS.n320 45.6589
R11541 VSS.n369 VSS.n368 44.4317
R11542 VSS.n368 VSS.n367 44.4317
R11543 VSS.n366 VSS.n365 44.4317
R11544 VSS.n365 VSS.n364 44.4317
R11545 VSS.n364 VSS.n363 44.4317
R11546 VSS.n363 VSS.n362 44.4317
R11547 VSS.n362 VSS.n361 44.4317
R11548 VSS.n361 VSS.t17 44.4317
R11549 VSS.n2900 VSS.n2899 44.4317
R11550 VSS.n2901 VSS.n2900 44.4317
R11551 VSS.n2902 VSS.n2901 44.4317
R11552 VSS.n2903 VSS.n2902 44.4317
R11553 VSS.n2904 VSS.n2903 44.4317
R11554 VSS.n2906 VSS.n2905 44.4317
R11555 VSS.n2907 VSS.n2906 44.4317
R11556 VSS.n2268 VSS.n2263 39.5975
R11557 VSS.n373 VSS.n358 39.2828
R11558 VSS.n367 VSS.t15 37.8977
R11559 VSS.n2905 VSS.t23 37.8977
R11560 VSS.n47 VSS.n46 35.3887
R11561 VSS.n70 VSS.n69 34.6307
R11562 VSS.n810 VSS.n808 33.0932
R11563 VSS.n823 VSS.n822 32.781
R11564 VSS.n2914 VSS.n2897 32.6533
R11565 VSS.n990 VSS.n988 32.3053
R11566 VSS.n1001 VSS.n1000 32.3053
R11567 VSS.n1121 VSS.n1119 32.3053
R11568 VSS.n1132 VSS.n1131 32.3053
R11569 VSS.n1224 VSS.n1222 32.3053
R11570 VSS.n1235 VSS.n1234 32.3053
R11571 VSS.n1347 VSS.n1345 32.3053
R11572 VSS.n1358 VSS.n1357 32.3053
R11573 VSS.n1478 VSS.n1477 32.3053
R11574 VSS.n671 VSS.n669 32.3053
R11575 VSS.n682 VSS.n681 32.3053
R11576 VSS.n22 VSS.n21 32.3053
R11577 VSS.n1593 VSS.n1592 32.3053
R11578 VSS.n358 VSS.n356 32.2375
R11579 VSS.n356 VSS.n354 32.2375
R11580 VSS.n354 VSS.n352 32.2375
R11581 VSS.n352 VSS.n350 32.2375
R11582 VSS.n350 VSS.n348 32.2375
R11583 VSS.n348 VSS.n346 32.2375
R11584 VSS.n346 VSS.n344 32.2375
R11585 VSS.n344 VSS.n342 32.2375
R11586 VSS.n342 VSS.n340 32.2375
R11587 VSS.n2249 VSS.n2247 32.2375
R11588 VSS.n2251 VSS.n2249 32.2375
R11589 VSS.n2253 VSS.n2251 32.2375
R11590 VSS.n2255 VSS.n2253 32.2375
R11591 VSS.n2257 VSS.n2255 32.2375
R11592 VSS.n2259 VSS.n2257 32.2375
R11593 VSS.n2261 VSS.n2259 32.2375
R11594 VSS.n2263 VSS.n2261 32.2375
R11595 VSS.n149 VSS.n147 31.8066
R11596 VSS.n523 VSS.n521 31.554
R11597 VSS.n222 VSS.n221 31.554
R11598 VSS.n536 VSS.n535 31.2563
R11599 VSS.n147 VSS.n145 26.3763
R11600 VSS.n145 VSS.n143 26.3763
R11601 VSS.n143 VSS.n141 26.3763
R11602 VSS.n141 VSS.n139 26.3763
R11603 VSS.n139 VSS.n137 26.3763
R11604 VSS.n137 VSS.n135 26.3763
R11605 VSS.n135 VSS.n133 26.3763
R11606 VSS.n133 VSS.n131 26.3763
R11607 VSS.n131 VSS.n129 26.3763
R11608 VSS.n2883 VSS.n2881 26.3763
R11609 VSS.n2885 VSS.n2883 26.3763
R11610 VSS.n2887 VSS.n2885 26.3763
R11611 VSS.n2889 VSS.n2887 26.3763
R11612 VSS.n2891 VSS.n2889 26.3763
R11613 VSS.n2893 VSS.n2891 26.3763
R11614 VSS.n2895 VSS.n2893 26.3763
R11615 VSS.n2897 VSS.n2895 26.3763
R11616 VSS.n1452 VSS.t8 23.4155
R11617 VSS.n1101 VSS.t13 23.4133
R11618 VSS.n654 VSS.t3 23.0658
R11619 VSS.n654 VSS.t4 23.0531
R11620 VSS.n68 VSS.t5 21.5627
R11621 VSS.n2908 VSS.t0 21.5627
R11622 VSS.n3359 VSS.t2 21.5627
R11623 VSS.n812 VSS.n810 21.2298
R11624 VSS.n814 VSS.n812 21.2298
R11625 VSS.n818 VSS.n814 21.2298
R11626 VSS.n820 VSS.n818 21.2298
R11627 VSS.n822 VSS.n820 21.2298
R11628 VSS.n39 VSS.n38 20.9093
R11629 VSS.n992 VSS.n990 20.7243
R11630 VSS.n994 VSS.n992 20.7243
R11631 VSS.n996 VSS.n994 20.7243
R11632 VSS.n998 VSS.n996 20.7243
R11633 VSS.n1000 VSS.n998 20.7243
R11634 VSS.n1123 VSS.n1121 20.7243
R11635 VSS.n1125 VSS.n1123 20.7243
R11636 VSS.n1127 VSS.n1125 20.7243
R11637 VSS.n1129 VSS.n1127 20.7243
R11638 VSS.n1131 VSS.n1129 20.7243
R11639 VSS.n1226 VSS.n1224 20.7243
R11640 VSS.n1228 VSS.n1226 20.7243
R11641 VSS.n1230 VSS.n1228 20.7243
R11642 VSS.n1232 VSS.n1230 20.7243
R11643 VSS.n1234 VSS.n1232 20.7243
R11644 VSS.n1349 VSS.n1347 20.7243
R11645 VSS.n1351 VSS.n1349 20.7243
R11646 VSS.n1353 VSS.n1351 20.7243
R11647 VSS.n1355 VSS.n1353 20.7243
R11648 VSS.n1357 VSS.n1355 20.7243
R11649 VSS.n1469 VSS.n1467 20.7243
R11650 VSS.n1471 VSS.n1469 20.7243
R11651 VSS.n1473 VSS.n1471 20.7243
R11652 VSS.n1475 VSS.n1473 20.7243
R11653 VSS.n1477 VSS.n1475 20.7243
R11654 VSS.n673 VSS.n671 20.7243
R11655 VSS.n675 VSS.n673 20.7243
R11656 VSS.n677 VSS.n675 20.7243
R11657 VSS.n679 VSS.n677 20.7243
R11658 VSS.n681 VSS.n679 20.7243
R11659 VSS.n1586 VSS.n1584 20.7243
R11660 VSS.n1588 VSS.n1586 20.7243
R11661 VSS.n1590 VSS.n1588 20.7243
R11662 VSS.n1592 VSS.n1590 20.7243
R11663 VSS.n525 VSS.n523 20.2424
R11664 VSS.n527 VSS.n525 20.2424
R11665 VSS.n531 VSS.n527 20.2424
R11666 VSS.n533 VSS.n531 20.2424
R11667 VSS.n535 VSS.n533 20.2424
R11668 VSS.n213 VSS.n211 20.2424
R11669 VSS.n215 VSS.n213 20.2424
R11670 VSS.n217 VSS.n215 20.2424
R11671 VSS.n219 VSS.n217 20.2424
R11672 VSS.n221 VSS.n219 20.2424
R11673 VSS.n312 VSS.n309 19.0364
R11674 VSS.n309 VSS.n308 18.8723
R11675 VSS.n669 VSS.n663 18.8723
R11676 VSS.n669 VSS.n668 18.8723
R11677 VSS.n988 VSS.n982 18.8723
R11678 VSS.n988 VSS.n987 18.8723
R11679 VSS.n1119 VSS.n1112 18.8723
R11680 VSS.n1119 VSS.n1118 18.8723
R11681 VSS.n1222 VSS.n1216 18.8723
R11682 VSS.n1222 VSS.n1221 18.8723
R11683 VSS.n1345 VSS.n1341 18.8723
R11684 VSS.n1345 VSS.n1344 18.8723
R11685 VSS.n8 VSS.n7 18.8723
R11686 VSS.n11 VSS.n8 18.8723
R11687 VSS.n22 VSS.n19 18.8723
R11688 VSS.n25 VSS.n22 18.8723
R11689 VSS.n808 VSS.n807 18.6666
R11690 VSS.n521 VSS.n520 18.4714
R11691 VSS.n808 VSS.n802 18.4714
R11692 VSS.n1878 VSS.t51 16.5305
R11693 VSS.n1878 VSS.t43 16.5305
R11694 VSS.n1869 VSS.t135 16.5305
R11695 VSS.n1869 VSS.t91 16.5305
R11696 VSS.n1860 VSS.t70 16.5305
R11697 VSS.n1860 VSS.t62 16.5305
R11698 VSS.n1851 VSS.t16 16.5305
R11699 VSS.n1851 VSS.t114 16.5305
R11700 VSS.n1842 VSS.t107 16.5305
R11701 VSS.n1842 VSS.t65 16.5305
R11702 VSS.n1833 VSS.t36 16.5305
R11703 VSS.n1833 VSS.t118 16.5305
R11704 VSS.n1824 VSS.t109 16.5305
R11705 VSS.n1824 VSS.t81 16.5305
R11706 VSS.n1815 VSS.t40 16.5305
R11707 VSS.n1815 VSS.t28 16.5305
R11708 VSS.n1806 VSS.t87 16.5305
R11709 VSS.n1806 VSS.t83 16.5305
R11710 VSS.n1797 VSS.t88 16.5305
R11711 VSS.n1797 VSS.t53 16.5305
R11712 VSS.n1788 VSS.t19 16.5305
R11713 VSS.n1788 VSS.t98 16.5305
R11714 VSS.n1779 VSS.t110 16.5305
R11715 VSS.n1779 VSS.t25 16.5305
R11716 VSS.n1770 VSS.t132 16.5305
R11717 VSS.n1770 VSS.t123 16.5305
R11718 VSS.n1761 VSS.t86 16.5305
R11719 VSS.n1761 VSS.t93 16.5305
R11720 VSS.n1752 VSS.t131 16.5305
R11721 VSS.n1752 VSS.t136 16.5305
R11722 VSS.n1743 VSS.t27 16.5305
R11723 VSS.n1743 VSS.t78 16.5305
R11724 VSS.n1734 VSS.t89 16.5305
R11725 VSS.n1734 VSS.t55 16.5305
R11726 VSS.n1725 VSS.t42 16.5305
R11727 VSS.n1725 VSS.t84 16.5305
R11728 VSS.n1716 VSS.t112 16.5305
R11729 VSS.n1716 VSS.t29 16.5305
R11730 VSS.n1707 VSS.t39 16.5305
R11731 VSS.n1707 VSS.t48 16.5305
R11732 VSS.n195 VSS.t138 16.5305
R11733 VSS.n182 VSS.t12 16.5305
R11734 VSS.n169 VSS.t9 16.5305
R11735 VSS.n169 VSS.t7 16.5305
R11736 VSS.n156 VSS.t6 16.5305
R11737 VSS.n2057 VSS.t117 16.5305
R11738 VSS.n2057 VSS.t106 16.5305
R11739 VSS.n2048 VSS.t74 16.5305
R11740 VSS.n2048 VSS.t35 16.5305
R11741 VSS.n2039 VSS.t130 16.5305
R11742 VSS.n2039 VSS.t127 16.5305
R11743 VSS.n2030 VSS.t82 16.5305
R11744 VSS.n2030 VSS.t59 16.5305
R11745 VSS.n2021 VSS.t52 16.5305
R11746 VSS.n2021 VSS.t129 16.5305
R11747 VSS.n2012 VSS.t99 16.5305
R11748 VSS.n2012 VSS.t60 16.5305
R11749 VSS.n2003 VSS.t56 16.5305
R11750 VSS.n2003 VSS.t20 16.5305
R11751 VSS.n1994 VSS.t102 16.5305
R11752 VSS.n1994 VSS.t96 16.5305
R11753 VSS.n1985 VSS.t30 16.5305
R11754 VSS.n1985 VSS.t21 16.5305
R11755 VSS.n1976 VSS.t32 16.5305
R11756 VSS.n1976 VSS.t120 16.5305
R11757 VSS.n1967 VSS.t85 16.5305
R11758 VSS.n1967 VSS.t44 16.5305
R11759 VSS.n1958 VSS.t57 16.5305
R11760 VSS.n1958 VSS.t92 16.5305
R11761 VSS.n1949 VSS.t73 16.5305
R11762 VSS.n1949 VSS.t63 16.5305
R11763 VSS.n1940 VSS.t26 16.5305
R11764 VSS.n1940 VSS.t38 16.5305
R11765 VSS.n1931 VSS.t72 16.5305
R11766 VSS.n1931 VSS.t75 16.5305
R11767 VSS.n1922 VSS.t95 16.5305
R11768 VSS.n1922 VSS.t18 16.5305
R11769 VSS.n1913 VSS.t33 16.5305
R11770 VSS.n1913 VSS.t122 16.5305
R11771 VSS.n1904 VSS.t103 16.5305
R11772 VSS.n1904 VSS.t22 16.5305
R11773 VSS.n1895 VSS.t58 16.5305
R11774 VSS.n1895 VSS.t97 16.5305
R11775 VSS.n1886 VSS.t101 16.5305
R11776 VSS.n1886 VSS.t111 16.5305
R11777 VSS.n2236 VSS.t125 16.5305
R11778 VSS.n2236 VSS.t121 16.5305
R11779 VSS.n2227 VSS.t79 16.5305
R11780 VSS.n2227 VSS.t49 16.5305
R11781 VSS.n2218 VSS.t137 16.5305
R11782 VSS.n2218 VSS.t133 16.5305
R11783 VSS.n2209 VSS.t90 16.5305
R11784 VSS.n2209 VSS.t68 16.5305
R11785 VSS.n2200 VSS.t61 16.5305
R11786 VSS.n2200 VSS.t134 16.5305
R11787 VSS.n2191 VSS.t113 16.5305
R11788 VSS.n2191 VSS.t69 16.5305
R11789 VSS.n2182 VSS.t64 16.5305
R11790 VSS.n2182 VSS.t31 16.5305
R11791 VSS.n2173 VSS.t116 16.5305
R11792 VSS.n2173 VSS.t105 16.5305
R11793 VSS.n2164 VSS.t45 16.5305
R11794 VSS.n2164 VSS.t34 16.5305
R11795 VSS.n2155 VSS.t46 16.5305
R11796 VSS.n2155 VSS.t126 16.5305
R11797 VSS.n2146 VSS.t94 16.5305
R11798 VSS.n2146 VSS.t54 16.5305
R11799 VSS.n2137 VSS.t66 16.5305
R11800 VSS.n2137 VSS.t100 16.5305
R11801 VSS.n2128 VSS.t77 16.5305
R11802 VSS.n2128 VSS.t71 16.5305
R11803 VSS.n2119 VSS.t41 16.5305
R11804 VSS.n2119 VSS.t50 16.5305
R11805 VSS.n2110 VSS.t76 16.5305
R11806 VSS.n2110 VSS.t80 16.5305
R11807 VSS.n2101 VSS.t104 16.5305
R11808 VSS.n2101 VSS.t24 16.5305
R11809 VSS.n2092 VSS.t47 16.5305
R11810 VSS.n2092 VSS.t128 16.5305
R11811 VSS.n2083 VSS.t119 16.5305
R11812 VSS.n2083 VSS.t37 16.5305
R11813 VSS.n2074 VSS.t67 16.5305
R11814 VSS.n2074 VSS.t108 16.5305
R11815 VSS.n2065 VSS.t115 16.5305
R11816 VSS.n2065 VSS.t124 16.5305
R11817 VSS.n44 VSS.n36 16.3383
R11818 VSS.n65 VSS.t11 15.0287
R11819 VSS.t1 VSS.n67 15.0287
R11820 VSS.n1879 VSS.n1878 11.6553
R11821 VSS.n1870 VSS.n1869 11.6553
R11822 VSS.n1861 VSS.n1860 11.6553
R11823 VSS.n1852 VSS.n1851 11.6553
R11824 VSS.n1843 VSS.n1842 11.6553
R11825 VSS.n1834 VSS.n1833 11.6553
R11826 VSS.n1825 VSS.n1824 11.6553
R11827 VSS.n1816 VSS.n1815 11.6553
R11828 VSS.n1807 VSS.n1806 11.6553
R11829 VSS.n1798 VSS.n1797 11.6553
R11830 VSS.n1789 VSS.n1788 11.6553
R11831 VSS.n1780 VSS.n1779 11.6553
R11832 VSS.n1771 VSS.n1770 11.6553
R11833 VSS.n1762 VSS.n1761 11.6553
R11834 VSS.n1753 VSS.n1752 11.6553
R11835 VSS.n1744 VSS.n1743 11.6553
R11836 VSS.n1735 VSS.n1734 11.6553
R11837 VSS.n1726 VSS.n1725 11.6553
R11838 VSS.n1717 VSS.n1716 11.6553
R11839 VSS.n1708 VSS.n1707 11.6553
R11840 VSS.n2058 VSS.n2057 11.6553
R11841 VSS.n2049 VSS.n2048 11.6553
R11842 VSS.n2040 VSS.n2039 11.6553
R11843 VSS.n2031 VSS.n2030 11.6553
R11844 VSS.n2022 VSS.n2021 11.6553
R11845 VSS.n2013 VSS.n2012 11.6553
R11846 VSS.n2004 VSS.n2003 11.6553
R11847 VSS.n1995 VSS.n1994 11.6553
R11848 VSS.n1986 VSS.n1985 11.6553
R11849 VSS.n1977 VSS.n1976 11.6553
R11850 VSS.n1968 VSS.n1967 11.6553
R11851 VSS.n1959 VSS.n1958 11.6553
R11852 VSS.n1950 VSS.n1949 11.6553
R11853 VSS.n1941 VSS.n1940 11.6553
R11854 VSS.n1932 VSS.n1931 11.6553
R11855 VSS.n1923 VSS.n1922 11.6553
R11856 VSS.n1914 VSS.n1913 11.6553
R11857 VSS.n1905 VSS.n1904 11.6553
R11858 VSS.n1896 VSS.n1895 11.6553
R11859 VSS.n1887 VSS.n1886 11.6553
R11860 VSS.n2237 VSS.n2236 11.6553
R11861 VSS.n2228 VSS.n2227 11.6553
R11862 VSS.n2219 VSS.n2218 11.6553
R11863 VSS.n2210 VSS.n2209 11.6553
R11864 VSS.n2201 VSS.n2200 11.6553
R11865 VSS.n2192 VSS.n2191 11.6553
R11866 VSS.n2183 VSS.n2182 11.6553
R11867 VSS.n2174 VSS.n2173 11.6553
R11868 VSS.n2165 VSS.n2164 11.6553
R11869 VSS.n2156 VSS.n2155 11.6553
R11870 VSS.n2147 VSS.n2146 11.6553
R11871 VSS.n2138 VSS.n2137 11.6553
R11872 VSS.n2129 VSS.n2128 11.6553
R11873 VSS.n2120 VSS.n2119 11.6553
R11874 VSS.n2111 VSS.n2110 11.6553
R11875 VSS.n2102 VSS.n2101 11.6553
R11876 VSS.n2093 VSS.n2092 11.6553
R11877 VSS.n2084 VSS.n2083 11.6553
R11878 VSS.n2075 VSS.n2074 11.6553
R11879 VSS.n2066 VSS.n2065 11.6553
R11880 VSS.n43 VSS.n42 11.2946
R11881 VSS.n320 VSS.n317 11.1595
R11882 VSS.n317 VSS.n315 11.1595
R11883 VSS.n315 VSS.n312 11.1595
R11884 VSS.n308 VSS.n305 11.1595
R11885 VSS.n305 VSS.n302 11.1595
R11886 VSS.n302 VSS.n300 11.1595
R11887 VSS.n807 VSS.n804 11.1595
R11888 VSS.n663 VSS.n659 11.1595
R11889 VSS.n668 VSS.n665 11.1595
R11890 VSS.n982 VSS.n978 11.1595
R11891 VSS.n987 VSS.n984 11.1595
R11892 VSS.n1112 VSS.n1109 11.1595
R11893 VSS.n1118 VSS.n1114 11.1595
R11894 VSS.n1216 VSS.n1212 11.1595
R11895 VSS.n1221 VSS.n1218 11.1595
R11896 VSS.n1341 VSS.n1338 11.1595
R11897 VSS.n4 VSS.n2 11.1595
R11898 VSS.n7 VSS.n4 11.1595
R11899 VSS.n14 VSS.n11 11.1595
R11900 VSS.n16 VSS.n14 11.1595
R11901 VSS.n19 VSS.n16 11.1595
R11902 VSS.n28 VSS.n25 11.1595
R11903 VSS.n30 VSS.n28 11.1595
R11904 VSS.n36 VSS.n30 11.1595
R11905 VSS.n520 VSS.n517 11.0182
R11906 VSS.n517 VSS.n515 11.0182
R11907 VSS.n515 VSS.n512 11.0182
R11908 VSS.n512 VSS.n509 11.0182
R11909 VSS.n509 VSS.n507 11.0182
R11910 VSS.n794 VSS.n792 11.0182
R11911 VSS.n797 VSS.n794 11.0182
R11912 VSS.n799 VSS.n797 11.0182
R11913 VSS.n802 VSS.n799 11.0182
R11914 VSS.n198 VSS.n197 9.3005
R11915 VSS.n185 VSS.n184 9.3005
R11916 VSS.n172 VSS.n171 9.3005
R11917 VSS.n159 VSS.n158 9.3005
R11918 VSS.n72 VSS.n70 9.14811
R11919 VSS.n157 VSS.n156 8.77119
R11920 VSS.n170 VSS.n169 8.63765
R11921 VSS.n196 VSS.n195 8.49781
R11922 VSS.n183 VSS.n182 8.49781
R11923 VSS.n44 VSS.n43 7.85619
R11924 VSS.n2274 VSS.n2273 7.82508
R11925 VSS.n3421 VSS.t14 7.18791
R11926 VSS.n3396 VSS.t10 7.18791
R11927 VSS.n67 VSS.n66 6.53451
R11928 VSS.t15 VSS.n366 6.53451
R11929 VSS.t23 VSS.n2904 6.53451
R11930 VSS.n333 VSS.n332 5.74009
R11931 VSS.n3369 VSS.n3368 5.5968
R11932 VSS.n153 VSS.n127 4.93165
R11933 VSS.n2926 VSS.n2922 4.73086
R11934 VSS.n2879 VSS.n2878 4.6505
R11935 VSS.n2875 VSS.n2874 4.6505
R11936 VSS.n2868 VSS.n2867 4.6505
R11937 VSS.n2861 VSS.n2860 4.6505
R11938 VSS.n2854 VSS.n2853 4.6505
R11939 VSS.n2847 VSS.n2846 4.6505
R11940 VSS.n2840 VSS.n2839 4.6505
R11941 VSS.n2832 VSS.n2831 4.6505
R11942 VSS.n2826 VSS.n2825 4.6505
R11943 VSS.n2816 VSS.n2815 4.6505
R11944 VSS.n2810 VSS.n2809 4.6505
R11945 VSS.n2802 VSS.n2801 4.6505
R11946 VSS.n2796 VSS.n2795 4.6505
R11947 VSS.n2788 VSS.n2787 4.6505
R11948 VSS.n2782 VSS.n2781 4.6505
R11949 VSS.n2772 VSS.n2771 4.6505
R11950 VSS.n2766 VSS.n2765 4.6505
R11951 VSS.n2758 VSS.n2757 4.6505
R11952 VSS.n2751 VSS.n2750 4.6505
R11953 VSS.n2744 VSS.n2743 4.6505
R11954 VSS.n2737 VSS.n2736 4.6505
R11955 VSS.n2730 VSS.n2729 4.6505
R11956 VSS.n2723 VSS.n2722 4.6505
R11957 VSS.n2716 VSS.n2715 4.6505
R11958 VSS.n2708 VSS.n2707 4.6505
R11959 VSS.n2702 VSS.n2701 4.6505
R11960 VSS.n2692 VSS.n2691 4.6505
R11961 VSS.n2686 VSS.n2685 4.6505
R11962 VSS.n2678 VSS.n2677 4.6505
R11963 VSS.n2672 VSS.n2671 4.6505
R11964 VSS.n2664 VSS.n2663 4.6505
R11965 VSS.n2658 VSS.n2657 4.6505
R11966 VSS.n2648 VSS.n2647 4.6505
R11967 VSS.n2642 VSS.n2641 4.6505
R11968 VSS.n2634 VSS.n2633 4.6505
R11969 VSS.n2627 VSS.n2626 4.6505
R11970 VSS.n2620 VSS.n2619 4.6505
R11971 VSS.n2613 VSS.n2612 4.6505
R11972 VSS.n2606 VSS.n2605 4.6505
R11973 VSS.n2599 VSS.n2598 4.6505
R11974 VSS.n2592 VSS.n2591 4.6505
R11975 VSS.n2584 VSS.n2583 4.6505
R11976 VSS.n2578 VSS.n2577 4.6505
R11977 VSS.n2568 VSS.n2567 4.6505
R11978 VSS.n2562 VSS.n2561 4.6505
R11979 VSS.n2554 VSS.n2553 4.6505
R11980 VSS.n2548 VSS.n2547 4.6505
R11981 VSS.n2540 VSS.n2539 4.6505
R11982 VSS.n2534 VSS.n2533 4.6505
R11983 VSS.n2524 VSS.n2523 4.6505
R11984 VSS.n2518 VSS.n2517 4.6505
R11985 VSS.n2510 VSS.n2509 4.6505
R11986 VSS.n2503 VSS.n2502 4.6505
R11987 VSS.n2496 VSS.n2495 4.6505
R11988 VSS.n2489 VSS.n2488 4.6505
R11989 VSS.n2482 VSS.n2481 4.6505
R11990 VSS.n2475 VSS.n2474 4.6505
R11991 VSS.n2468 VSS.n2467 4.6505
R11992 VSS.n2460 VSS.n2459 4.6505
R11993 VSS.n2454 VSS.n2453 4.6505
R11994 VSS.n2444 VSS.n2443 4.6505
R11995 VSS.n2438 VSS.n2437 4.6505
R11996 VSS.n2430 VSS.n2429 4.6505
R11997 VSS.n2424 VSS.n2423 4.6505
R11998 VSS.n2416 VSS.n2415 4.6505
R11999 VSS.n2410 VSS.n2409 4.6505
R12000 VSS.n2400 VSS.n2399 4.6505
R12001 VSS.n2394 VSS.n2393 4.6505
R12002 VSS.n2386 VSS.n2385 4.6505
R12003 VSS.n2379 VSS.n2378 4.6505
R12004 VSS.n2372 VSS.n2371 4.6505
R12005 VSS.n2365 VSS.n2364 4.6505
R12006 VSS.n2358 VSS.n2357 4.6505
R12007 VSS.n2351 VSS.n2350 4.6505
R12008 VSS.n2344 VSS.n2343 4.6505
R12009 VSS.n2336 VSS.n2335 4.6505
R12010 VSS.n2330 VSS.n2329 4.6505
R12011 VSS.n2320 VSS.n2319 4.6505
R12012 VSS.n2314 VSS.n2313 4.6505
R12013 VSS.n2306 VSS.n2305 4.6505
R12014 VSS.n2300 VSS.n2299 4.6505
R12015 VSS.n2292 VSS.n2291 4.6505
R12016 VSS.n2286 VSS.n2285 4.6505
R12017 VSS.n2276 VSS.n2275 4.6505
R12018 VSS.n2975 VSS.n2974 4.6505
R12019 VSS.n2973 VSS.n2972 4.6505
R12020 VSS.n2969 VSS.n2968 4.6505
R12021 VSS.n2965 VSS.n2964 4.6505
R12022 VSS.n2961 VSS.n2960 4.6505
R12023 VSS.n2957 VSS.n2956 4.6505
R12024 VSS.n2953 VSS.n2952 4.6505
R12025 VSS.n2949 VSS.n2948 4.6505
R12026 VSS.n2945 VSS.n2944 4.6505
R12027 VSS.n2938 VSS.n2937 4.6505
R12028 VSS.n2934 VSS.n2933 4.6505
R12029 VSS.n2930 VSS.n2929 4.6505
R12030 VSS.n2926 VSS.n2925 4.6505
R12031 VSS.n2981 VSS.n2980 4.6505
R12032 VSS.n2986 VSS.n2985 4.6505
R12033 VSS.n2990 VSS.n2989 4.6505
R12034 VSS.n2995 VSS.n2994 4.6505
R12035 VSS.n3000 VSS.n2999 4.6505
R12036 VSS.n3004 VSS.n3003 4.6505
R12037 VSS.n3009 VSS.n3008 4.6505
R12038 VSS.n3015 VSS.n3014 4.6505
R12039 VSS.n3020 VSS.n3019 4.6505
R12040 VSS.n3024 VSS.n3023 4.6505
R12041 VSS.n3029 VSS.n3028 4.6505
R12042 VSS.n3033 VSS.n3032 4.6505
R12043 VSS.n3038 VSS.n3037 4.6505
R12044 VSS.n3042 VSS.n3041 4.6505
R12045 VSS.n3047 VSS.n3046 4.6505
R12046 VSS.n3052 VSS.n3051 4.6505
R12047 VSS.n3056 VSS.n3055 4.6505
R12048 VSS.n3061 VSS.n3060 4.6505
R12049 VSS.n3065 VSS.n3064 4.6505
R12050 VSS.n3070 VSS.n3069 4.6505
R12051 VSS.n3074 VSS.n3073 4.6505
R12052 VSS.n3079 VSS.n3078 4.6505
R12053 VSS.n3083 VSS.n3082 4.6505
R12054 VSS.n3088 VSS.n3087 4.6505
R12055 VSS.n3094 VSS.n3093 4.6505
R12056 VSS.n3099 VSS.n3098 4.6505
R12057 VSS.n3103 VSS.n3102 4.6505
R12058 VSS.n3108 VSS.n3107 4.6505
R12059 VSS.n3112 VSS.n3111 4.6505
R12060 VSS.n3117 VSS.n3116 4.6505
R12061 VSS.n3121 VSS.n3120 4.6505
R12062 VSS.n3126 VSS.n3125 4.6505
R12063 VSS.n3131 VSS.n3130 4.6505
R12064 VSS.n3135 VSS.n3134 4.6505
R12065 VSS.n3140 VSS.n3139 4.6505
R12066 VSS.n3144 VSS.n3143 4.6505
R12067 VSS.n3149 VSS.n3148 4.6505
R12068 VSS.n3153 VSS.n3152 4.6505
R12069 VSS.n3158 VSS.n3157 4.6505
R12070 VSS.n3162 VSS.n3161 4.6505
R12071 VSS.n3167 VSS.n3166 4.6505
R12072 VSS.n3173 VSS.n3172 4.6505
R12073 VSS.n3178 VSS.n3177 4.6505
R12074 VSS.n3182 VSS.n3181 4.6505
R12075 VSS.n3187 VSS.n3186 4.6505
R12076 VSS.n3191 VSS.n3190 4.6505
R12077 VSS.n3196 VSS.n3195 4.6505
R12078 VSS.n3200 VSS.n3199 4.6505
R12079 VSS.n3205 VSS.n3204 4.6505
R12080 VSS.n3210 VSS.n3209 4.6505
R12081 VSS.n3214 VSS.n3213 4.6505
R12082 VSS.n3219 VSS.n3218 4.6505
R12083 VSS.n3223 VSS.n3222 4.6505
R12084 VSS.n3228 VSS.n3227 4.6505
R12085 VSS.n3232 VSS.n3231 4.6505
R12086 VSS.n3237 VSS.n3236 4.6505
R12087 VSS.n3241 VSS.n3240 4.6505
R12088 VSS.n3246 VSS.n3245 4.6505
R12089 VSS.n3252 VSS.n3251 4.6505
R12090 VSS.n3257 VSS.n3256 4.6505
R12091 VSS.n3261 VSS.n3260 4.6505
R12092 VSS.n3266 VSS.n3265 4.6505
R12093 VSS.n3270 VSS.n3269 4.6505
R12094 VSS.n3275 VSS.n3274 4.6505
R12095 VSS.n3279 VSS.n3278 4.6505
R12096 VSS.n3284 VSS.n3283 4.6505
R12097 VSS.n3289 VSS.n3288 4.6505
R12098 VSS.n3293 VSS.n3292 4.6505
R12099 VSS.n3298 VSS.n3297 4.6505
R12100 VSS.n3302 VSS.n3301 4.6505
R12101 VSS.n3307 VSS.n3306 4.6505
R12102 VSS.n3311 VSS.n3310 4.6505
R12103 VSS.n3316 VSS.n3315 4.6505
R12104 VSS.n3320 VSS.n3319 4.6505
R12105 VSS.n3325 VSS.n3324 4.6505
R12106 VSS.n3331 VSS.n3330 4.6505
R12107 VSS.n3336 VSS.n3335 4.6505
R12108 VSS.n3340 VSS.n3339 4.6505
R12109 VSS.n3345 VSS.n3344 4.6505
R12110 VSS.n3349 VSS.n3348 4.6505
R12111 VSS.n3354 VSS.n3353 4.6505
R12112 VSS.n3358 VSS.n3357 4.6505
R12113 VSS.n3365 VSS.n3364 4.6505
R12114 VSS.n3367 VSS.n3366 4.6505
R12115 VSS.n2917 VSS.n2916 4.6505
R12116 VSS.n3440 VSS.n3439 4.6505
R12117 VSS.n3435 VSS.n3434 4.6505
R12118 VSS.n3430 VSS.n3429 4.6505
R12119 VSS.n3425 VSS.n3424 4.6505
R12120 VSS.n3420 VSS.n3419 4.6505
R12121 VSS.n3415 VSS.n3414 4.6505
R12122 VSS.n3410 VSS.n3409 4.6505
R12123 VSS.n3405 VSS.n3404 4.6505
R12124 VSS.n3400 VSS.n3399 4.6505
R12125 VSS.n3395 VSS.n3394 4.6505
R12126 VSS.n3390 VSS.n3389 4.6505
R12127 VSS.n3385 VSS.n3384 4.6505
R12128 VSS.n3380 VSS.n3379 4.6505
R12129 VSS.n3375 VSS.n3374 4.6505
R12130 VSS.n3371 VSS.n3370 4.6505
R12131 VSS.n3449 VSS.n3448 4.6505
R12132 VSS.n2919 VSS.n2918 4.6505
R12133 VSS.n3445 VSS.n3444 4.6505
R12134 VSS.n691 VSS.n656 4.51047
R12135 VSS.n1712 VSS.n1711 4.5005
R12136 VSS.n1721 VSS.n1720 4.5005
R12137 VSS.n1730 VSS.n1729 4.5005
R12138 VSS.n1739 VSS.n1738 4.5005
R12139 VSS.n1748 VSS.n1747 4.5005
R12140 VSS.n1757 VSS.n1756 4.5005
R12141 VSS.n1766 VSS.n1765 4.5005
R12142 VSS.n1775 VSS.n1774 4.5005
R12143 VSS.n1784 VSS.n1783 4.5005
R12144 VSS.n1793 VSS.n1792 4.5005
R12145 VSS.n1802 VSS.n1801 4.5005
R12146 VSS.n1811 VSS.n1810 4.5005
R12147 VSS.n1820 VSS.n1819 4.5005
R12148 VSS.n1829 VSS.n1828 4.5005
R12149 VSS.n1838 VSS.n1837 4.5005
R12150 VSS.n1847 VSS.n1846 4.5005
R12151 VSS.n1856 VSS.n1855 4.5005
R12152 VSS.n1865 VSS.n1864 4.5005
R12153 VSS.n1874 VSS.n1873 4.5005
R12154 VSS.n1883 VSS.n1882 4.5005
R12155 VSS.n202 VSS.n201 4.5005
R12156 VSS.n189 VSS.n188 4.5005
R12157 VSS.n176 VSS.n175 4.5005
R12158 VSS.n163 VSS.n162 4.5005
R12159 VSS.n1663 VSS.n1662 4.5005
R12160 VSS.n1658 VSS.n1657 4.5005
R12161 VSS.n1648 VSS.n1647 4.5005
R12162 VSS.n1635 VSS.n1634 4.5005
R12163 VSS.n1599 VSS.n1598 4.5005
R12164 VSS.n1578 VSS.n1577 4.5005
R12165 VSS.n1568 VSS.n1567 4.5005
R12166 VSS.n1525 VSS.n1524 4.5005
R12167 VSS.n1533 VSS.n1532 4.5005
R12168 VSS.n1517 VSS.n1516 4.5005
R12169 VSS.n1507 VSS.n1506 4.5005
R12170 VSS.n1494 VSS.n1493 4.5005
R12171 VSS.n1450 VSS.n1449 4.5005
R12172 VSS.n1439 VSS.n1438 4.5005
R12173 VSS.n1426 VSS.n1425 4.5005
R12174 VSS.n1384 VSS.n1383 4.5005
R12175 VSS.n1389 VSS.n1388 4.5005
R12176 VSS.n1373 VSS.n1372 4.5005
R12177 VSS.n1364 VSS.n1363 4.5005
R12178 VSS.n1332 VSS.n1331 4.5005
R12179 VSS.n1300 VSS.n1299 4.5005
R12180 VSS.n1286 VSS.n1285 4.5005
R12181 VSS.n1274 VSS.n1273 4.5005
R12182 VSS.n1208 VSS.n1207 4.5005
R12183 VSS.n1241 VSS.n1240 4.5005
R12184 VSS.n1203 VSS.n1202 4.5005
R12185 VSS.n1194 VSS.n1193 4.5005
R12186 VSS.n1179 VSS.n1178 4.5005
R12187 VSS.n1147 VSS.n1146 4.5005
R12188 VSS.n1136 VSS.n1135 4.5005
R12189 VSS.n1100 VSS.n1099 4.5005
R12190 VSS.n1057 VSS.n1056 4.5005
R12191 VSS.n1065 VSS.n1064 4.5005
R12192 VSS.n1049 VSS.n1048 4.5005
R12193 VSS.n1037 VSS.n1036 4.5005
R12194 VSS.n1024 VSS.n1023 4.5005
R12195 VSS.n970 VSS.n969 4.5005
R12196 VSS.n957 VSS.n956 4.5005
R12197 VSS.n945 VSS.n944 4.5005
R12198 VSS.n903 VSS.n902 4.5005
R12199 VSS.n911 VSS.n910 4.5005
R12200 VSS.n896 VSS.n895 4.5005
R12201 VSS.n691 VSS.n690 4.5005
R12202 VSS.n864 VSS.n863 4.5005
R12203 VSS.n851 VSS.n850 4.5005
R12204 VSS.n838 VSS.n837 4.5005
R12205 VSS.n827 VSS.n826 4.5005
R12206 VSS.n831 VSS.n830 4.5005
R12207 VSS.n787 VSS.n786 4.5005
R12208 VSS.n777 VSS.n776 4.5005
R12209 VSS.n764 VSS.n763 4.5005
R12210 VSS.n731 VSS.n730 4.5005
R12211 VSS.n717 VSS.n716 4.5005
R12212 VSS.n705 VSS.n704 4.5005
R12213 VSS.n593 VSS.n592 4.5005
R12214 VSS.n697 VSS.n696 4.5005
R12215 VSS.n586 VSS.n585 4.5005
R12216 VSS.n577 VSS.n576 4.5005
R12217 VSS.n563 VSS.n562 4.5005
R12218 VSS.n502 VSS.n501 4.5005
R12219 VSS.n491 VSS.n490 4.5005
R12220 VSS.n477 VSS.n476 4.5005
R12221 VSS.n434 VSS.n433 4.5005
R12222 VSS.n439 VSS.n438 4.5005
R12223 VSS.n423 VSS.n422 4.5005
R12224 VSS.n416 VSS.n415 4.5005
R12225 VSS.n228 VSS.n227 4.5005
R12226 VSS.n262 VSS.n261 4.5005
R12227 VSS.n275 VSS.n274 4.5005
R12228 VSS.n284 VSS.n283 4.5005
R12229 VSS.n1891 VSS.n1890 4.5005
R12230 VSS.n1900 VSS.n1899 4.5005
R12231 VSS.n1909 VSS.n1908 4.5005
R12232 VSS.n1918 VSS.n1917 4.5005
R12233 VSS.n1927 VSS.n1926 4.5005
R12234 VSS.n1936 VSS.n1935 4.5005
R12235 VSS.n1945 VSS.n1944 4.5005
R12236 VSS.n1954 VSS.n1953 4.5005
R12237 VSS.n1963 VSS.n1962 4.5005
R12238 VSS.n1972 VSS.n1971 4.5005
R12239 VSS.n1981 VSS.n1980 4.5005
R12240 VSS.n1990 VSS.n1989 4.5005
R12241 VSS.n1999 VSS.n1998 4.5005
R12242 VSS.n2008 VSS.n2007 4.5005
R12243 VSS.n2017 VSS.n2016 4.5005
R12244 VSS.n2026 VSS.n2025 4.5005
R12245 VSS.n2035 VSS.n2034 4.5005
R12246 VSS.n2044 VSS.n2043 4.5005
R12247 VSS.n2053 VSS.n2052 4.5005
R12248 VSS.n2062 VSS.n2061 4.5005
R12249 VSS.n2070 VSS.n2069 4.5005
R12250 VSS.n2079 VSS.n2078 4.5005
R12251 VSS.n2088 VSS.n2087 4.5005
R12252 VSS.n2097 VSS.n2096 4.5005
R12253 VSS.n2106 VSS.n2105 4.5005
R12254 VSS.n2115 VSS.n2114 4.5005
R12255 VSS.n2124 VSS.n2123 4.5005
R12256 VSS.n2133 VSS.n2132 4.5005
R12257 VSS.n2142 VSS.n2141 4.5005
R12258 VSS.n2151 VSS.n2150 4.5005
R12259 VSS.n2160 VSS.n2159 4.5005
R12260 VSS.n2169 VSS.n2168 4.5005
R12261 VSS.n2178 VSS.n2177 4.5005
R12262 VSS.n2187 VSS.n2186 4.5005
R12263 VSS.n2196 VSS.n2195 4.5005
R12264 VSS.n2205 VSS.n2204 4.5005
R12265 VSS.n2214 VSS.n2213 4.5005
R12266 VSS.n2223 VSS.n2222 4.5005
R12267 VSS.n2232 VSS.n2231 4.5005
R12268 VSS.n2241 VSS.n2240 4.5005
R12269 VSS.n529 VSS.n528 3.89846
R12270 VSS.n816 VSS.n815 3.7456
R12271 VSS.n2915 VSS.n2914 3.73591
R12272 VSS.n3014 VSS.n3011 3.73383
R12273 VSS.n3093 VSS.n3090 3.73383
R12274 VSS.n3172 VSS.n3169 3.73383
R12275 VSS.n3251 VSS.n3248 3.73383
R12276 VSS.n3330 VSS.n3327 3.73383
R12277 VSS.n3014 VSS.n3013 3.5205
R12278 VSS.n3093 VSS.n3092 3.5205
R12279 VSS.n3172 VSS.n3171 3.5205
R12280 VSS.n3251 VSS.n3250 3.5205
R12281 VSS.n3330 VSS.n3329 3.5205
R12282 VSS.n3008 VSS.n3007 3.30717
R12283 VSS.n3087 VSS.n3086 3.30717
R12284 VSS.n3166 VSS.n3165 3.30717
R12285 VSS.n3245 VSS.n3244 3.30717
R12286 VSS.n3324 VSS.n3323 3.30717
R12287 VSS.n2269 VSS.n2268 3.18987
R12288 VSS.n2979 VSS.n2978 3.10915
R12289 VSS.n3019 VSS.n3018 3.09383
R12290 VSS.n3098 VSS.n3097 3.09383
R12291 VSS.n3177 VSS.n3176 3.09383
R12292 VSS.n3256 VSS.n3255 3.09383
R12293 VSS.n3335 VSS.n3334 3.09383
R12294 VSS.n1626 VSS.n1625 3.03311
R12295 VSS.n1610 VSS.n1609 3.03311
R12296 VSS.n1483 VSS.n1482 3.03311
R12297 VSS.n1461 VSS.n1460 3.03311
R12298 VSS.n1325 VSS.n1324 3.03311
R12299 VSS.n1310 VSS.n1309 3.03311
R12300 VSS.n1169 VSS.n1168 3.03311
R12301 VSS.n1157 VSS.n1156 3.03311
R12302 VSS.n1014 VSS.n1013 3.03311
R12303 VSS.n1003 VSS.n1002 3.03311
R12304 VSS.n886 VSS.n885 3.03311
R12305 VSS.n875 VSS.n874 3.03311
R12306 VSS.n755 VSS.n754 3.03311
R12307 VSS.n741 VSS.n740 3.03311
R12308 VSS.n552 VSS.n551 3.03311
R12309 VSS.n540 VSS.n539 3.03311
R12310 VSS.n238 VSS.n237 3.03311
R12311 VSS.n251 VSS.n250 3.03311
R12312 VSS.n691 VSS.n687 3.02303
R12313 VSS.n1882 VSS.n1881 3.01226
R12314 VSS.n1873 VSS.n1872 3.01226
R12315 VSS.n1864 VSS.n1863 3.01226
R12316 VSS.n1855 VSS.n1854 3.01226
R12317 VSS.n1846 VSS.n1845 3.01226
R12318 VSS.n1837 VSS.n1836 3.01226
R12319 VSS.n1828 VSS.n1827 3.01226
R12320 VSS.n1819 VSS.n1818 3.01226
R12321 VSS.n1810 VSS.n1809 3.01226
R12322 VSS.n1801 VSS.n1800 3.01226
R12323 VSS.n1792 VSS.n1791 3.01226
R12324 VSS.n1783 VSS.n1782 3.01226
R12325 VSS.n1774 VSS.n1773 3.01226
R12326 VSS.n1765 VSS.n1764 3.01226
R12327 VSS.n1756 VSS.n1755 3.01226
R12328 VSS.n1747 VSS.n1746 3.01226
R12329 VSS.n1738 VSS.n1737 3.01226
R12330 VSS.n1729 VSS.n1728 3.01226
R12331 VSS.n1720 VSS.n1719 3.01226
R12332 VSS.n1711 VSS.n1710 3.01226
R12333 VSS.n2061 VSS.n2060 3.01226
R12334 VSS.n2052 VSS.n2051 3.01226
R12335 VSS.n2043 VSS.n2042 3.01226
R12336 VSS.n2034 VSS.n2033 3.01226
R12337 VSS.n2025 VSS.n2024 3.01226
R12338 VSS.n2016 VSS.n2015 3.01226
R12339 VSS.n2007 VSS.n2006 3.01226
R12340 VSS.n1998 VSS.n1997 3.01226
R12341 VSS.n1989 VSS.n1988 3.01226
R12342 VSS.n1980 VSS.n1979 3.01226
R12343 VSS.n1971 VSS.n1970 3.01226
R12344 VSS.n1962 VSS.n1961 3.01226
R12345 VSS.n1953 VSS.n1952 3.01226
R12346 VSS.n1944 VSS.n1943 3.01226
R12347 VSS.n1935 VSS.n1934 3.01226
R12348 VSS.n1926 VSS.n1925 3.01226
R12349 VSS.n1917 VSS.n1916 3.01226
R12350 VSS.n1908 VSS.n1907 3.01226
R12351 VSS.n1899 VSS.n1898 3.01226
R12352 VSS.n1890 VSS.n1889 3.01226
R12353 VSS.n2240 VSS.n2239 3.01226
R12354 VSS.n2231 VSS.n2230 3.01226
R12355 VSS.n2222 VSS.n2221 3.01226
R12356 VSS.n2213 VSS.n2212 3.01226
R12357 VSS.n2204 VSS.n2203 3.01226
R12358 VSS.n2195 VSS.n2194 3.01226
R12359 VSS.n2186 VSS.n2185 3.01226
R12360 VSS.n2177 VSS.n2176 3.01226
R12361 VSS.n2168 VSS.n2167 3.01226
R12362 VSS.n2159 VSS.n2158 3.01226
R12363 VSS.n2150 VSS.n2149 3.01226
R12364 VSS.n2141 VSS.n2140 3.01226
R12365 VSS.n2132 VSS.n2131 3.01226
R12366 VSS.n2123 VSS.n2122 3.01226
R12367 VSS.n2114 VSS.n2113 3.01226
R12368 VSS.n2105 VSS.n2104 3.01226
R12369 VSS.n2096 VSS.n2095 3.01226
R12370 VSS.n2087 VSS.n2086 3.01226
R12371 VSS.n2078 VSS.n2077 3.01226
R12372 VSS.n2069 VSS.n2068 3.01226
R12373 VSS.n2273 VSS.n2271 2.89219
R12374 VSS.n3003 VSS.n3002 2.8805
R12375 VSS.n3082 VSS.n3081 2.8805
R12376 VSS.n3161 VSS.n3160 2.8805
R12377 VSS.n3240 VSS.n3239 2.8805
R12378 VSS.n3319 VSS.n3318 2.8805
R12379 VSS.n47 VSS.n44 2.8677
R12380 VSS.n152 VSS.n149 2.66944
R12381 VSS.n3023 VSS.n3022 2.66717
R12382 VSS.n3102 VSS.n3101 2.66717
R12383 VSS.n3181 VSS.n3180 2.66717
R12384 VSS.n3260 VSS.n3259 2.66717
R12385 VSS.n3339 VSS.n3338 2.66717
R12386 VSS.n2999 VSS.n2998 2.45383
R12387 VSS.n3078 VSS.n3077 2.45383
R12388 VSS.n3157 VSS.n3156 2.45383
R12389 VSS.n3236 VSS.n3235 2.45383
R12390 VSS.n3315 VSS.n3314 2.45383
R12391 VSS.n1460 VSS.n1456 2.41559
R12392 VSS.n2329 VSS.n2322 2.36572
R12393 VSS.n2453 VSS.n2446 2.36572
R12394 VSS.n2577 VSS.n2571 2.36572
R12395 VSS.n2701 VSS.n2695 2.36572
R12396 VSS.n2825 VSS.n2819 2.36572
R12397 VSS.n53 VSS.n49 2.32157
R12398 VSS.n191 VSS.n183 2.30562
R12399 VSS.n204 VSS.n196 2.30538
R12400 VSS.n2285 VSS.n2284 2.29615
R12401 VSS.n2409 VSS.n2408 2.29615
R12402 VSS.n2533 VSS.n2532 2.29615
R12403 VSS.n2657 VSS.n2656 2.29615
R12404 VSS.n2781 VSS.n2780 2.29615
R12405 VSS.n178 VSS.n170 2.26697
R12406 VSS.n3028 VSS.n3027 2.2405
R12407 VSS.n3107 VSS.n3106 2.2405
R12408 VSS.n3186 VSS.n3185 2.2405
R12409 VSS.n3265 VSS.n3264 2.2405
R12410 VSS.n3344 VSS.n3343 2.2405
R12411 VSS.n165 VSS.n157 2.22907
R12412 VSS.n1324 VSS.n1323 2.22239
R12413 VSS.n2319 VSS.n2316 2.08746
R12414 VSS.n2443 VSS.n2440 2.08746
R12415 VSS.n2567 VSS.n2564 2.08746
R12416 VSS.n2691 VSS.n2688 2.08746
R12417 VSS.n2815 VSS.n2812 2.08746
R12418 VSS.n1013 VSS.n1012 2.02918
R12419 VSS.n2994 VSS.n2993 2.02717
R12420 VSS.n3073 VSS.n3072 2.02717
R12421 VSS.n3152 VSS.n3151 2.02717
R12422 VSS.n3231 VSS.n3230 2.02717
R12423 VSS.n3310 VSS.n3309 2.02717
R12424 VSS.n2291 VSS.n2290 2.01789
R12425 VSS.n2415 VSS.n2414 2.01789
R12426 VSS.n2539 VSS.n2538 2.01789
R12427 VSS.n2663 VSS.n2662 2.01789
R12428 VSS.n2787 VSS.n2786 2.01789
R12429 VSS.n58 VSS.n56 1.9461
R12430 VSS.n62 VSS.n60 1.9461
R12431 VSS.n374 VSS.n373 1.94572
R12432 VSS.n296 VSS.n295 1.93258
R12433 VSS.n96 VSS.n94 1.85241
R12434 VSS.n120 VSS.n117 1.85241
R12435 VSS.n122 VSS.n120 1.85241
R12436 VSS.n754 VSS.n753 1.84292
R12437 VSS.n1624 VSS.n1619 1.83597
R12438 VSS.n3032 VSS.n3031 1.81383
R12439 VSS.n3111 VSS.n3110 1.81383
R12440 VSS.n3190 VSS.n3189 1.81383
R12441 VSS.n3269 VSS.n3268 1.81383
R12442 VSS.n3348 VSS.n3347 1.81383
R12443 VSS.n2313 VSS.n2309 1.8092
R12444 VSS.n2437 VSS.n2433 1.8092
R12445 VSS.n2561 VSS.n2557 1.8092
R12446 VSS.n2685 VSS.n2681 1.8092
R12447 VSS.n2809 VSS.n2805 1.8092
R12448 VSS.n127 VSS.n125 1.78411
R12449 VSS.n125 VSS.n124 1.77833
R12450 VSS.n2281 VSS.n2278 1.73963
R12451 VSS.n2299 VSS.n2298 1.73963
R12452 VSS.n2328 VSS.n2325 1.73963
R12453 VSS.n2334 VSS.n2332 1.73963
R12454 VSS.n2342 VSS.n2339 1.73963
R12455 VSS.n2392 VSS.n2389 1.73963
R12456 VSS.n2398 VSS.n2396 1.73963
R12457 VSS.n2405 VSS.n2402 1.73963
R12458 VSS.n2423 VSS.n2422 1.73963
R12459 VSS.n2452 VSS.n2449 1.73963
R12460 VSS.n2458 VSS.n2456 1.73963
R12461 VSS.n2466 VSS.n2463 1.73963
R12462 VSS.n2516 VSS.n2513 1.73963
R12463 VSS.n2522 VSS.n2520 1.73963
R12464 VSS.n2529 VSS.n2526 1.73963
R12465 VSS.n2547 VSS.n2546 1.73963
R12466 VSS.n2576 VSS.n2573 1.73963
R12467 VSS.n2582 VSS.n2580 1.73963
R12468 VSS.n2590 VSS.n2587 1.73963
R12469 VSS.n2640 VSS.n2637 1.73963
R12470 VSS.n2646 VSS.n2644 1.73963
R12471 VSS.n2653 VSS.n2650 1.73963
R12472 VSS.n2671 VSS.n2670 1.73963
R12473 VSS.n2700 VSS.n2697 1.73963
R12474 VSS.n2706 VSS.n2704 1.73963
R12475 VSS.n2714 VSS.n2711 1.73963
R12476 VSS.n2764 VSS.n2761 1.73963
R12477 VSS.n2770 VSS.n2768 1.73963
R12478 VSS.n2777 VSS.n2774 1.73963
R12479 VSS.n2795 VSS.n2794 1.73963
R12480 VSS.n2824 VSS.n2821 1.73963
R12481 VSS.n2830 VSS.n2828 1.73963
R12482 VSS.n2838 VSS.n2835 1.73963
R12483 VSS.n3448 VSS.n3447 1.69389
R12484 VSS.n1002 VSS.n1001 1.69107
R12485 VSS.n237 VSS.n233 1.64276
R12486 VSS.n237 VSS.n236 1.64276
R12487 VSS.n2276 VSS.n2274 1.64141
R12488 VSS.n330 VSS.n328 1.63352
R12489 VSS.n324 VSS.n322 1.63352
R12490 VSS.n326 VSS.n324 1.63352
R12491 VSS.n328 VSS.n326 1.63352
R12492 VSS.n332 VSS.n330 1.63352
R12493 VSS.n154 VSS.n122 1.60731
R12494 VSS.n2385 VSS.n2381 1.6005
R12495 VSS.n2509 VSS.n2505 1.6005
R12496 VSS.n2633 VSS.n2629 1.6005
R12497 VSS.n2757 VSS.n2753 1.6005
R12498 VSS.n2878 VSS.n2877 1.6005
R12499 VSS.n786 VSS.n784 1.6005
R12500 VSS.n2989 VSS.n2988 1.6005
R12501 VSS.n3069 VSS.n3068 1.6005
R12502 VSS.n3148 VSS.n3147 1.6005
R12503 VSS.n3227 VSS.n3226 1.6005
R12504 VSS.n3306 VSS.n3305 1.6005
R12505 VSS.n2305 VSS.n2302 1.53093
R12506 VSS.n2350 VSS.n2349 1.53093
R12507 VSS.n2429 VSS.n2426 1.53093
R12508 VSS.n2474 VSS.n2473 1.53093
R12509 VSS.n2553 VSS.n2550 1.53093
R12510 VSS.n2598 VSS.n2597 1.53093
R12511 VSS.n2677 VSS.n2674 1.53093
R12512 VSS.n2722 VSS.n2721 1.53093
R12513 VSS.n2801 VSS.n2798 1.53093
R12514 VSS.n2846 VSS.n2845 1.53093
R12515 VSS.n1697 VSS.n1696 1.5005
R12516 VSS.n1704 VSS.n1703 1.5005
R12517 VSS.n3444 VSS.n3443 1.49466
R12518 VSS.n2305 VSS.n2304 1.46137
R12519 VSS.n2429 VSS.n2428 1.46137
R12520 VSS.n2553 VSS.n2552 1.46137
R12521 VSS.n2677 VSS.n2676 1.46137
R12522 VSS.n2801 VSS.n2800 1.46137
R12523 VSS.n250 VSS.n245 1.44956
R12524 VSS.n2944 VSS.n2941 1.44635
R12525 VSS.n1036 VSS.n1030 1.40125
R12526 VSS.n1048 VSS.n1044 1.40125
R12527 VSS.n1482 VSS.n1478 1.40125
R12528 VSS.n3037 VSS.n3036 1.38717
R12529 VSS.n3116 VSS.n3115 1.38717
R12530 VSS.n3195 VSS.n3194 1.38717
R12531 VSS.n3274 VSS.n3273 1.38717
R12532 VSS.n3353 VSS.n3352 1.38717
R12533 VSS.n100 VSS.n97 1.3622
R12534 VSS.n2937 VSS.n2936 1.3613
R12535 VSS.n2944 VSS.n2943 1.3613
R12536 VSS.n550 VSS.n547 1.35808
R12537 VSS.n750 VSS.n747 1.35808
R12538 VSS.n773 VSS.n770 1.35808
R12539 VSS.n115 VSS.n112 1.33497
R12540 VSS.n2378 VSS.n2375 1.32224
R12541 VSS.n2502 VSS.n2499 1.32224
R12542 VSS.n2626 VSS.n2623 1.32224
R12543 VSS.n2750 VSS.n2747 1.32224
R12544 VSS.n2874 VSS.n2871 1.32224
R12545 VSS.n3439 VSS.n3438 1.29544
R12546 VSS.n3374 VSS.n3373 1.29544
R12547 VSS.n740 VSS.n737 1.26111
R12548 VSS.n1013 VSS.n1010 1.25635
R12549 VSS.n104 VSS.n101 1.25327
R12550 VSS.n2299 VSS.n2295 1.25267
R12551 VSS.n2357 VSS.n2356 1.25267
R12552 VSS.n2423 VSS.n2419 1.25267
R12553 VSS.n2481 VSS.n2480 1.25267
R12554 VSS.n2547 VSS.n2543 1.25267
R12555 VSS.n2605 VSS.n2604 1.25267
R12556 VSS.n2671 VSS.n2667 1.25267
R12557 VSS.n2729 VSS.n2728 1.25267
R12558 VSS.n2795 VSS.n2791 1.25267
R12559 VSS.n2853 VSS.n2852 1.25267
R12560 VSS.n1363 VSS.n1360 1.20805
R12561 VSS.n1372 VSS.n1370 1.20805
R12562 VSS.n2933 VSS.n2932 1.1912
R12563 VSS.n2948 VSS.n2947 1.1912
R12564 VSS.n2313 VSS.n2312 1.18311
R12565 VSS.n2437 VSS.n2436 1.18311
R12566 VSS.n2561 VSS.n2560 1.18311
R12567 VSS.n2685 VSS.n2684 1.18311
R12568 VSS.n2809 VSS.n2808 1.18311
R12569 VSS.n2985 VSS.n2984 1.17383
R12570 VSS.n3064 VSS.n3063 1.17383
R12571 VSS.n3143 VSS.n3142 1.17383
R12572 VSS.n3222 VSS.n3221 1.17383
R12573 VSS.n3301 VSS.n3300 1.17383
R12574 VSS.n1884 VSS.n1883 1.13663
R12575 VSS.n1875 VSS.n1874 1.13663
R12576 VSS.n1866 VSS.n1865 1.13663
R12577 VSS.n1857 VSS.n1856 1.13663
R12578 VSS.n1848 VSS.n1847 1.13663
R12579 VSS.n1839 VSS.n1838 1.13663
R12580 VSS.n1830 VSS.n1829 1.13663
R12581 VSS.n1821 VSS.n1820 1.13663
R12582 VSS.n1812 VSS.n1811 1.13663
R12583 VSS.n1803 VSS.n1802 1.13663
R12584 VSS.n1794 VSS.n1793 1.13663
R12585 VSS.n1785 VSS.n1784 1.13663
R12586 VSS.n1776 VSS.n1775 1.13663
R12587 VSS.n1767 VSS.n1766 1.13663
R12588 VSS.n1758 VSS.n1757 1.13663
R12589 VSS.n1749 VSS.n1748 1.13663
R12590 VSS.n1740 VSS.n1739 1.13663
R12591 VSS.n1731 VSS.n1730 1.13663
R12592 VSS.n1722 VSS.n1721 1.13663
R12593 VSS.n1713 VSS.n1712 1.13663
R12594 VSS.n2063 VSS.n2062 1.13663
R12595 VSS.n2054 VSS.n2053 1.13663
R12596 VSS.n2045 VSS.n2044 1.13663
R12597 VSS.n2036 VSS.n2035 1.13663
R12598 VSS.n2027 VSS.n2026 1.13663
R12599 VSS.n2018 VSS.n2017 1.13663
R12600 VSS.n2009 VSS.n2008 1.13663
R12601 VSS.n2000 VSS.n1999 1.13663
R12602 VSS.n1991 VSS.n1990 1.13663
R12603 VSS.n1982 VSS.n1981 1.13663
R12604 VSS.n1973 VSS.n1972 1.13663
R12605 VSS.n1964 VSS.n1963 1.13663
R12606 VSS.n1955 VSS.n1954 1.13663
R12607 VSS.n1946 VSS.n1945 1.13663
R12608 VSS.n1937 VSS.n1936 1.13663
R12609 VSS.n1928 VSS.n1927 1.13663
R12610 VSS.n1919 VSS.n1918 1.13663
R12611 VSS.n1910 VSS.n1909 1.13663
R12612 VSS.n1901 VSS.n1900 1.13663
R12613 VSS.n1892 VSS.n1891 1.13663
R12614 VSS.n2242 VSS.n2241 1.13663
R12615 VSS.n2233 VSS.n2232 1.13663
R12616 VSS.n2224 VSS.n2223 1.13663
R12617 VSS.n2215 VSS.n2214 1.13663
R12618 VSS.n2206 VSS.n2205 1.13663
R12619 VSS.n2197 VSS.n2196 1.13663
R12620 VSS.n2188 VSS.n2187 1.13663
R12621 VSS.n2179 VSS.n2178 1.13663
R12622 VSS.n2170 VSS.n2169 1.13663
R12623 VSS.n2161 VSS.n2160 1.13663
R12624 VSS.n2152 VSS.n2151 1.13663
R12625 VSS.n2143 VSS.n2142 1.13663
R12626 VSS.n2134 VSS.n2133 1.13663
R12627 VSS.n2125 VSS.n2124 1.13663
R12628 VSS.n2116 VSS.n2115 1.13663
R12629 VSS.n2107 VSS.n2106 1.13663
R12630 VSS.n2098 VSS.n2097 1.13663
R12631 VSS.n2089 VSS.n2088 1.13663
R12632 VSS.n2080 VSS.n2079 1.13663
R12633 VSS.n2071 VSS.n2070 1.13663
R12634 VSS.n441 VSS.n440 1.1255
R12635 VSS.n595 VSS.n594 1.1255
R12636 VSS.n913 VSS.n912 1.1255
R12637 VSS.n1067 VSS.n1066 1.1255
R12638 VSS.n1243 VSS.n1242 1.1255
R12639 VSS.n1391 VSS.n1390 1.1255
R12640 VSS.n1535 VSS.n1534 1.1255
R12641 VSS.n1681 VSS.n1680 1.1255
R12642 VSS.n3434 VSS.n3433 1.09622
R12643 VSS.n3379 VSS.n3378 1.09622
R12644 VSS.n49 VSS.n47 1.09277
R12645 VSS.n1002 VSS.n976 1.06314
R12646 VSS.n2371 VSS.n2367 1.04398
R12647 VSS.n2495 VSS.n2491 1.04398
R12648 VSS.n2619 VSS.n2615 1.04398
R12649 VSS.n2743 VSS.n2739 1.04398
R12650 VSS.n2867 VSS.n2863 1.04398
R12651 VSS.n2929 VSS.n2928 1.0211
R12652 VSS.n2952 VSS.n2951 1.0211
R12653 VSS.n1647 VSS.n1641 1.01484
R12654 VSS.n1657 VSS.n1655 1.01484
R12655 VSS.n2291 VSS.n2288 0.974413
R12656 VSS.n2364 VSS.n2363 0.974413
R12657 VSS.n2415 VSS.n2412 0.974413
R12658 VSS.n2488 VSS.n2487 0.974413
R12659 VSS.n2539 VSS.n2536 0.974413
R12660 VSS.n2612 VSS.n2611 0.974413
R12661 VSS.n2663 VSS.n2660 0.974413
R12662 VSS.n2736 VSS.n2735 0.974413
R12663 VSS.n2787 VSS.n2784 0.974413
R12664 VSS.n2860 VSS.n2859 0.974413
R12665 VSS.n1240 VSS.n1235 0.966538
R12666 VSS.n1320 VSS.n1316 0.966538
R12667 VSS.n1383 VSS.n1382 0.966538
R12668 VSS.n1425 VSS.n1424 0.966538
R12669 VSS.n1438 VSS.n1437 0.966538
R12670 VSS.n3041 VSS.n3040 0.9605
R12671 VSS.n3120 VSS.n3119 0.9605
R12672 VSS.n3199 VSS.n3198 0.9605
R12673 VSS.n3278 VSS.n3277 0.9605
R12674 VSS.n3357 VSS.n3356 0.9605
R12675 VSS.n108 VSS.n62 0.9221
R12676 VSS.n2319 VSS.n2318 0.904848
R12677 VSS.n2443 VSS.n2442 0.904848
R12678 VSS.n2567 VSS.n2566 0.904848
R12679 VSS.n2691 VSS.n2690 0.904848
R12680 VSS.n2815 VSS.n2814 0.904848
R12681 VSS.n3429 VSS.n3428 0.896998
R12682 VSS.n3384 VSS.n3383 0.896998
R12683 VSS.n1309 VSS.n1306 0.869934
R12684 VSS.n1460 VSS.n1459 0.869934
R12685 VSS.n1625 VSS.n1617 0.869934
R12686 VSS.n2925 VSS.n2924 0.850998
R12687 VSS.n2956 VSS.n2955 0.850998
R12688 VSS.n683 VSS.n682 0.821632
R12689 VSS.n374 VSS.n333 0.81701
R12690 VSS.n205 VSS.n204 0.802347
R12691 VSS.n192 VSS.n191 0.802041
R12692 VSS.n179 VSS.n178 0.800604
R12693 VSS.n166 VSS.n165 0.79886
R12694 VSS.n561 VSS.n560 0.776258
R12695 VSS.n762 VSS.n761 0.776258
R12696 VSS.n226 VSS.n225 0.77333
R12697 VSS.n1056 VSS.n1055 0.77333
R12698 VSS.n1099 VSS.n1098 0.77333
R12699 VSS.n1135 VSS.n1134 0.77333
R12700 VSS.n1146 VSS.n1145 0.77333
R12701 VSS.n1330 VSS.n1329 0.77333
R12702 VSS.n1609 VSS.n1608 0.77333
R12703 VSS.n2978 VSS.n2977 0.765949
R12704 VSS.n2269 VSS.n2245 0.765717
R12705 VSS.n2364 VSS.n2361 0.765717
R12706 VSS.n2488 VSS.n2485 0.765717
R12707 VSS.n2612 VSS.n2609 0.765717
R12708 VSS.n2736 VSS.n2733 0.765717
R12709 VSS.n2860 VSS.n2857 0.765717
R12710 VSS.n3060 VSS.n3059 0.747167
R12711 VSS.n3139 VSS.n3138 0.747167
R12712 VSS.n3218 VSS.n3217 0.747167
R12713 VSS.n3297 VSS.n3296 0.747167
R12714 VSS.n86 VSS.n85 0.735819
R12715 VSS.n91 VSS.n90 0.735819
R12716 VSS.n726 VSS.n725 0.727773
R12717 VSS.n283 VSS.n282 0.725028
R12718 VSS.n274 VSS.n273 0.725028
R12719 VSS.n258 VSS.n257 0.725028
R12720 VSS.n261 VSS.n260 0.725028
R12721 VSS.n497 VSS.n496 0.725028
R12722 VSS.n1134 VSS.n1132 0.725028
R12723 VSS.n1142 VSS.n1141 0.725028
R12724 VSS.n1448 VSS.n1444 0.725028
R12725 VSS.n3424 VSS.n3423 0.697776
R12726 VSS.n3389 VSS.n3388 0.697776
R12727 VSS.n2285 VSS.n2281 0.696152
R12728 VSS.n2371 VSS.n2370 0.696152
R12729 VSS.n2409 VSS.n2405 0.696152
R12730 VSS.n2495 VSS.n2494 0.696152
R12731 VSS.n2533 VSS.n2529 0.696152
R12732 VSS.n2619 VSS.n2618 0.696152
R12733 VSS.n2657 VSS.n2653 0.696152
R12734 VSS.n2743 VSS.n2742 0.696152
R12735 VSS.n2781 VSS.n2777 0.696152
R12736 VSS.n2867 VSS.n2866 0.696152
R12737 VSS.n2922 VSS.n2921 0.680899
R12738 VSS.n2960 VSS.n2959 0.680899
R12739 VSS.n227 VSS.n222 0.676726
R12740 VSS.n225 VSS.n224 0.676726
R12741 VSS.n413 VSS.n412 0.676726
R12742 VSS.n686 VSS.n683 0.676726
R12743 VSS.n1295 VSS.n1294 0.676726
R12744 VSS.n1482 VSS.n1481 0.676726
R12745 VSS.n1609 VSS.n1605 0.676726
R12746 VSS.n85 VSS.n82 0.654117
R12747 VSS.n90 VSS.n88 0.654117
R12748 VSS.n105 VSS.n104 0.654117
R12749 VSS.n33 VSS.n32 0.653901
R12750 VSS.n38 VSS.n37 0.653901
R12751 VSS.n51 VSS.n50 0.653901
R12752 VSS.n66 VSS.n65 0.653901
R12753 VSS.t5 VSS.t1 0.653901
R12754 VSS.n69 VSS.n68 0.653901
R12755 VSS.n72 VSS.n71 0.653901
R12756 VSS.n75 VSS.n74 0.653901
R12757 VSS.n1621 VSS.n1620 0.653901
R12758 VSS.n250 VSS.n249 0.628425
R12759 VSS.n859 VSS.n856 0.628425
R12760 VSS.n2329 VSS.n2328 0.626587
R12761 VSS.n2453 VSS.n2452 0.626587
R12762 VSS.n2577 VSS.n2576 0.626587
R12763 VSS.n2701 VSS.n2700 0.626587
R12764 VSS.n2825 VSS.n2824 0.626587
R12765 VSS.n101 VSS.n100 0.599649
R12766 VSS.n2916 VSS.n2915 0.598165
R12767 VSS.n575 VSS.n574 0.582318
R12768 VSS.n775 VSS.n774 0.582318
R12769 VSS.n414 VSS.n413 0.580123
R12770 VSS.n539 VSS.n536 0.580123
R12771 VSS.n826 VSS.n825 0.580123
R12772 VSS.n837 VSS.n836 0.580123
R12773 VSS.n850 VSS.n849 0.580123
R12774 VSS.n863 VSS.n862 0.580123
R12775 VSS.n1362 VSS.n1361 0.580123
R12776 VSS.n1594 VSS.n1593 0.580123
R12777 VSS.n1625 VSS.n1624 0.580123
R12778 VSS.n375 VSS.n374 0.538425
R12779 VSS.n713 VSS.n712 0.533833
R12780 VSS.n3046 VSS.n3045 0.533833
R12781 VSS.n3125 VSS.n3124 0.533833
R12782 VSS.n3204 VSS.n3203 0.533833
R12783 VSS.n3283 VSS.n3282 0.533833
R12784 VSS.n3364 VSS.n3363 0.533833
R12785 VSS.n270 VSS.n269 0.531821
R12786 VSS.n271 VSS.n270 0.531821
R12787 VSS.n257 VSS.n256 0.531821
R12788 VSS.n483 VSS.n482 0.531821
R12789 VSS.n844 VSS.n843 0.531821
R12790 VSS.n1107 VSS.n1106 0.531821
R12791 VSS.n1432 VSS.n1431 0.531821
R12792 VSS.n112 VSS.n110 0.517947
R12793 VSS.n117 VSS.n115 0.517947
R12794 VSS.n2964 VSS.n2963 0.510799
R12795 VSS.n3419 VSS.n3418 0.498554
R12796 VSS.n3394 VSS.n3393 0.498554
R12797 VSS.n97 VSS.n96 0.490713
R12798 VSS.n2357 VSS.n2353 0.487457
R12799 VSS.n2481 VSS.n2477 0.487457
R12800 VSS.n2605 VSS.n2601 0.487457
R12801 VSS.n2729 VSS.n2725 0.487457
R12802 VSS.n2853 VSS.n2849 0.487457
R12803 VSS.n1880 VSS.n1879 0.487074
R12804 VSS.n1871 VSS.n1870 0.487074
R12805 VSS.n1862 VSS.n1861 0.487074
R12806 VSS.n1853 VSS.n1852 0.487074
R12807 VSS.n1844 VSS.n1843 0.487074
R12808 VSS.n1835 VSS.n1834 0.487074
R12809 VSS.n1826 VSS.n1825 0.487074
R12810 VSS.n1817 VSS.n1816 0.487074
R12811 VSS.n1808 VSS.n1807 0.487074
R12812 VSS.n1799 VSS.n1798 0.487074
R12813 VSS.n1790 VSS.n1789 0.487074
R12814 VSS.n1781 VSS.n1780 0.487074
R12815 VSS.n1772 VSS.n1771 0.487074
R12816 VSS.n1763 VSS.n1762 0.487074
R12817 VSS.n1754 VSS.n1753 0.487074
R12818 VSS.n1745 VSS.n1744 0.487074
R12819 VSS.n1736 VSS.n1735 0.487074
R12820 VSS.n1727 VSS.n1726 0.487074
R12821 VSS.n1718 VSS.n1717 0.487074
R12822 VSS.n1709 VSS.n1708 0.487074
R12823 VSS.n2059 VSS.n2058 0.487074
R12824 VSS.n2050 VSS.n2049 0.487074
R12825 VSS.n2041 VSS.n2040 0.487074
R12826 VSS.n2032 VSS.n2031 0.487074
R12827 VSS.n2023 VSS.n2022 0.487074
R12828 VSS.n2014 VSS.n2013 0.487074
R12829 VSS.n2005 VSS.n2004 0.487074
R12830 VSS.n1996 VSS.n1995 0.487074
R12831 VSS.n1987 VSS.n1986 0.487074
R12832 VSS.n1978 VSS.n1977 0.487074
R12833 VSS.n1969 VSS.n1968 0.487074
R12834 VSS.n1960 VSS.n1959 0.487074
R12835 VSS.n1951 VSS.n1950 0.487074
R12836 VSS.n1942 VSS.n1941 0.487074
R12837 VSS.n1933 VSS.n1932 0.487074
R12838 VSS.n1924 VSS.n1923 0.487074
R12839 VSS.n1915 VSS.n1914 0.487074
R12840 VSS.n1906 VSS.n1905 0.487074
R12841 VSS.n1897 VSS.n1896 0.487074
R12842 VSS.n1888 VSS.n1887 0.487074
R12843 VSS.n2238 VSS.n2237 0.487074
R12844 VSS.n2229 VSS.n2228 0.487074
R12845 VSS.n2220 VSS.n2219 0.487074
R12846 VSS.n2211 VSS.n2210 0.487074
R12847 VSS.n2202 VSS.n2201 0.487074
R12848 VSS.n2193 VSS.n2192 0.487074
R12849 VSS.n2184 VSS.n2183 0.487074
R12850 VSS.n2175 VSS.n2174 0.487074
R12851 VSS.n2166 VSS.n2165 0.487074
R12852 VSS.n2157 VSS.n2156 0.487074
R12853 VSS.n2148 VSS.n2147 0.487074
R12854 VSS.n2139 VSS.n2138 0.487074
R12855 VSS.n2130 VSS.n2129 0.487074
R12856 VSS.n2121 VSS.n2120 0.487074
R12857 VSS.n2112 VSS.n2111 0.487074
R12858 VSS.n2103 VSS.n2102 0.487074
R12859 VSS.n2094 VSS.n2093 0.487074
R12860 VSS.n2085 VSS.n2084 0.487074
R12861 VSS.n2076 VSS.n2075 0.487074
R12862 VSS.n2067 VSS.n2066 0.487074
R12863 VSS.n560 VSS.n559 0.485348
R12864 VSS.n574 VSS.n573 0.485348
R12865 VSS.n592 VSS.n589 0.485348
R12866 VSS.n704 VSS.n700 0.485348
R12867 VSS.n826 VSS.n790 0.4848
R12868 VSS.n297 VSS.n296 0.483519
R12869 VSS.n433 VSS.n426 0.483519
R12870 VSS.n476 VSS.n471 0.483519
R12871 VSS.n837 VSS.n834 0.483519
R12872 VSS.n874 VSS.n873 0.483519
R12873 VSS.n885 VSS.n882 0.483519
R12874 VSS.n902 VSS.n901 0.483519
R12875 VSS.n944 VSS.n943 0.483519
R12876 VSS.n1021 VSS.n1018 0.483519
R12877 VSS.n1034 VSS.n1031 0.483519
R12878 VSS.n1056 VSS.n1052 0.483519
R12879 VSS.n1099 VSS.n1096 0.483519
R12880 VSS.n1175 VSS.n1173 0.483519
R12881 VSS.n1187 VSS.n1184 0.483519
R12882 VSS.n1207 VSS.n1206 0.483519
R12883 VSS.n1273 VSS.n1272 0.483519
R12884 VSS.n1282 VSS.n1281 0.483519
R12885 VSS.n1492 VSS.n1491 0.483519
R12886 VSS.n1597 VSS.n1596 0.483519
R12887 VSS.n1662 VSS.n1661 0.483519
R12888 VSS.n404 VSS.n207 0.451649
R12889 VSS.n461 VSS.n194 0.450213
R12890 VSS.n601 VSS.n181 0.448776
R12891 VSS.n619 VSS.n168 0.447339
R12892 VSS.n585 VSS.n584 0.436864
R12893 VSS.n696 VSS.n695 0.436864
R12894 VSS.n786 VSS.n785 0.436864
R12895 VSS.n79 VSS.n78 0.436245
R12896 VSS.n149 VSS.n148 0.436245
R12897 VSS.n293 VSS.n292 0.435217
R12898 VSS.n422 VSS.n421 0.435217
R12899 VSS.n438 VSS.n437 0.435217
R12900 VSS.n830 VSS.n829 0.435217
R12901 VSS.n1372 VSS.n1371 0.435217
R12902 VSS.n1388 VSS.n1387 0.435217
R12903 VSS.n1516 VSS.n1515 0.435217
R12904 VSS.n1532 VSS.n1531 0.435217
R12905 VSS.n1657 VSS.n1656 0.435217
R12906 VSS.n155 VSS.n108 0.427322
R12907 VSS.n2378 VSS.n2377 0.417891
R12908 VSS.n2399 VSS.n2398 0.417891
R12909 VSS.n2502 VSS.n2501 0.417891
R12910 VSS.n2523 VSS.n2522 0.417891
R12911 VSS.n2626 VSS.n2625 0.417891
R12912 VSS.n2647 VSS.n2646 0.417891
R12913 VSS.n2750 VSS.n2749 0.417891
R12914 VSS.n2771 VSS.n2770 0.417891
R12915 VSS.n2874 VSS.n2873 0.417891
R12916 VSS.n3454 VSS.n1705 0.387366
R12917 VSS.n433 VSS.n432 0.386915
R12918 VSS.n476 VSS.n475 0.386915
R12919 VSS.n490 VSS.n489 0.386915
R12920 VSS.n501 VSS.n500 0.386915
R12921 VSS.n968 VSS.n967 0.386915
R12922 VSS.n1156 VSS.n1155 0.386915
R12923 VSS.n1379 VSS.n1376 0.386915
R12924 VSS.n1422 VSS.n1420 0.386915
R12925 VSS.n1524 VSS.n1523 0.386915
R12926 VSS.n1567 VSS.n1566 0.386915
R12927 VSS.n1633 VSS.n1632 0.386915
R12928 VSS.n1632 VSS.n1630 0.386915
R12929 VSS.n1645 VSS.n1642 0.386915
R12930 VSS.n201 VSS.n200 0.376971
R12931 VSS.n188 VSS.n187 0.376971
R12932 VSS.n175 VSS.n174 0.376971
R12933 VSS.n162 VSS.n161 0.376971
R12934 VSS.n56 VSS.n53 0.375967
R12935 VSS.n60 VSS.n58 0.375967
R12936 VSS.n107 VSS.n91 0.354543
R12937 VSS.n2335 VSS.n2334 0.348326
R12938 VSS.n2459 VSS.n2458 0.348326
R12939 VSS.n2583 VSS.n2582 0.348326
R12940 VSS.n2707 VSS.n2706 0.348326
R12941 VSS.n2831 VSS.n2830 0.348326
R12942 VSS.n108 VSS.n107 0.341833
R12943 VSS.n2968 VSS.n2967 0.340699
R12944 VSS.n712 VSS.n711 0.339894
R12945 VSS.n725 VSS.n724 0.339894
R12946 VSS.n954 VSS.n952 0.338613
R12947 VSS.n967 VSS.n964 0.338613
R12948 VSS.n1048 VSS.n1047 0.338613
R12949 VSS.n1064 VSS.n1063 0.338613
R12950 VSS.n1202 VSS.n1201 0.338613
R12951 VSS.n1240 VSS.n1239 0.338613
R12952 VSS.n3055 VSS.n3054 0.3205
R12953 VSS.n3134 VSS.n3133 0.3205
R12954 VSS.n3213 VSS.n3212 0.3205
R12955 VSS.n3292 VSS.n3291 0.3205
R12956 VSS.n655 VSS.n654 0.3005
R12957 VSS.n87 VSS.n86 0.300074
R12958 VSS.n3414 VSS.n3413 0.299333
R12959 VSS.n3399 VSS.n3398 0.299333
R12960 VSS.n716 VSS.n713 0.291409
R12961 VSS.n274 VSS.n271 0.290311
R12962 VSS.n490 VSS.n483 0.290311
R12963 VSS.n539 VSS.n538 0.290311
R12964 VSS.n825 VSS.n823 0.290311
R12965 VSS.n874 VSS.n870 0.290311
R12966 VSS.n885 VSS.n884 0.290311
R12967 VSS.n894 VSS.n891 0.290311
R12968 VSS.n909 VSS.n906 0.290311
R12969 VSS.n956 VSS.n955 0.290311
R12970 VSS.n1022 VSS.n1021 0.290311
R12971 VSS.n1135 VSS.n1107 0.290311
R12972 VSS.n1155 VSS.n1152 0.290311
R12973 VSS.n1167 VSS.n1164 0.290311
R12974 VSS.n1177 VSS.n1175 0.290311
R12975 VSS.n1285 VSS.n1282 0.290311
R12976 VSS.n1505 VSS.n1504 0.290311
R12977 VSS.n1576 VSS.n1575 0.290311
R12978 VSS.n1577 VSS.n1576 0.290311
R12979 VSS.n82 VSS.n81 0.27284
R12980 VSS.n376 VSS.n375 0.265654
R12981 VSS.n2274 VSS.n2269 0.25565
R12982 VSS.n80 VSS.n79 0.245606
R12983 VSS.n576 VSS.n575 0.242924
R12984 VSS.n763 VSS.n760 0.242924
R12985 VSS.n776 VSS.n773 0.242924
R12986 VSS.n776 VSS.n775 0.242924
R12987 VSS.n295 VSS.n293 0.242009
R12988 VSS.n415 VSS.n414 0.242009
R12989 VSS.n1036 VSS.n1035 0.242009
R12990 VSS.n1363 VSS.n1362 0.242009
R12991 VSS.n1506 VSS.n1505 0.242009
R12992 VSS.n1575 VSS.n1573 0.242009
R12993 VSS.n1596 VSS.n1594 0.242009
R12994 VSS.n1647 VSS.n1646 0.242009
R12995 VSS.n1714 VSS.n1713 0.227826
R12996 VSS.n1723 VSS.n1722 0.227826
R12997 VSS.n1732 VSS.n1731 0.227826
R12998 VSS.n1741 VSS.n1740 0.227826
R12999 VSS.n1750 VSS.n1749 0.227826
R13000 VSS.n1759 VSS.n1758 0.227826
R13001 VSS.n1768 VSS.n1767 0.227826
R13002 VSS.n1777 VSS.n1776 0.227826
R13003 VSS.n1786 VSS.n1785 0.227826
R13004 VSS.n1795 VSS.n1794 0.227826
R13005 VSS.n1804 VSS.n1803 0.227826
R13006 VSS.n1813 VSS.n1812 0.227826
R13007 VSS.n1822 VSS.n1821 0.227826
R13008 VSS.n1831 VSS.n1830 0.227826
R13009 VSS.n1840 VSS.n1839 0.227826
R13010 VSS.n1849 VSS.n1848 0.227826
R13011 VSS.n1858 VSS.n1857 0.227826
R13012 VSS.n1867 VSS.n1866 0.227826
R13013 VSS.n1876 VSS.n1875 0.227826
R13014 VSS.n1893 VSS.n1892 0.227826
R13015 VSS.n1902 VSS.n1901 0.227826
R13016 VSS.n1911 VSS.n1910 0.227826
R13017 VSS.n1920 VSS.n1919 0.227826
R13018 VSS.n1929 VSS.n1928 0.227826
R13019 VSS.n1938 VSS.n1937 0.227826
R13020 VSS.n1947 VSS.n1946 0.227826
R13021 VSS.n1956 VSS.n1955 0.227826
R13022 VSS.n1965 VSS.n1964 0.227826
R13023 VSS.n1974 VSS.n1973 0.227826
R13024 VSS.n1983 VSS.n1982 0.227826
R13025 VSS.n1992 VSS.n1991 0.227826
R13026 VSS.n2001 VSS.n2000 0.227826
R13027 VSS.n2010 VSS.n2009 0.227826
R13028 VSS.n2019 VSS.n2018 0.227826
R13029 VSS.n2028 VSS.n2027 0.227826
R13030 VSS.n2037 VSS.n2036 0.227826
R13031 VSS.n2046 VSS.n2045 0.227826
R13032 VSS.n2055 VSS.n2054 0.227826
R13033 VSS.n2072 VSS.n2071 0.227826
R13034 VSS.n2081 VSS.n2080 0.227826
R13035 VSS.n2090 VSS.n2089 0.227826
R13036 VSS.n2099 VSS.n2098 0.227826
R13037 VSS.n2108 VSS.n2107 0.227826
R13038 VSS.n2117 VSS.n2116 0.227826
R13039 VSS.n2126 VSS.n2125 0.227826
R13040 VSS.n2135 VSS.n2134 0.227826
R13041 VSS.n2144 VSS.n2143 0.227826
R13042 VSS.n2153 VSS.n2152 0.227826
R13043 VSS.n2162 VSS.n2161 0.227826
R13044 VSS.n2171 VSS.n2170 0.227826
R13045 VSS.n2180 VSS.n2179 0.227826
R13046 VSS.n2189 VSS.n2188 0.227826
R13047 VSS.n2198 VSS.n2197 0.227826
R13048 VSS.n2207 VSS.n2206 0.227826
R13049 VSS.n2216 VSS.n2215 0.227826
R13050 VSS.n2225 VSS.n2224 0.227826
R13051 VSS.n2234 VSS.n2233 0.227826
R13052 VSS.n153 VSS.n152 0.218372
R13053 VSS.n3453 VSS.n1884 0.216135
R13054 VSS.n3452 VSS.n2063 0.216135
R13055 VSS.n3451 VSS.n2242 0.216135
R13056 VSS.n3454 VSS.n3453 0.214983
R13057 VSS.n2350 VSS.n2347 0.209196
R13058 VSS.n2474 VSS.n2471 0.209196
R13059 VSS.n2598 VSS.n2595 0.209196
R13060 VSS.n2722 VSS.n2719 0.209196
R13061 VSS.n2846 VSS.n2843 0.209196
R13062 VSS.n592 VSS.n591 0.194439
R13063 VSS.n704 VSS.n703 0.194439
R13064 VSS.n716 VSS.n715 0.194439
R13065 VSS.n730 VSS.n729 0.194439
R13066 VSS.n292 VSS.n291 0.193708
R13067 VSS.n850 VSS.n846 0.193708
R13068 VSS.n955 VSS.n954 0.193708
R13069 VSS.n1168 VSS.n1167 0.193708
R13070 VSS.n1192 VSS.n1188 0.193708
R13071 VSS.n1285 VSS.n1284 0.193708
R13072 VSS.n1299 VSS.n1298 0.193708
R13073 VSS.n1434 VSS.n1432 0.193708
R13074 VSS.n1491 VSS.n1489 0.193708
R13075 VSS.n1504 VSS.n1502 0.193708
R13076 VSS.n1646 VSS.n1645 0.193708
R13077 VSS.n3453 VSS.n3452 0.193304
R13078 VSS.n3452 VSS.n3451 0.193304
R13079 VSS.n3451 VSS.n3450 0.173932
R13080 VSS.n2972 VSS.n2971 0.1706
R13081 VSS VSS.n155 0.169981
R13082 VSS.n88 VSS.n87 0.163904
R13083 VSS.n2979 VSS.n2976 0.160963
R13084 VSS.n2981 VSS.n2979 0.152767
R13085 VSS.n690 VSS.n689 0.145406
R13086 VSS.n895 VSS.n894 0.145406
R13087 VSS.n910 VSS.n909 0.145406
R13088 VSS.n952 VSS.n951 0.145406
R13089 VSS.n964 VSS.n963 0.145406
R13090 VSS.n2385 VSS.n2384 0.13963
R13091 VSS.n2393 VSS.n2392 0.13963
R13092 VSS.n2509 VSS.n2508 0.13963
R13093 VSS.n2517 VSS.n2516 0.13963
R13094 VSS.n2633 VSS.n2632 0.13963
R13095 VSS.n2641 VSS.n2640 0.13963
R13096 VSS.n2757 VSS.n2756 0.13963
R13097 VSS.n2765 VSS.n2764 0.13963
R13098 VSS.n78 VSS.n64 0.13667
R13099 VSS.n3371 VSS.n3369 0.130603
R13100 VSS.n687 VSS.n686 0.130042
R13101 VSS.n81 VSS.n80 0.109436
R13102 VSS.n3051 VSS.n3050 0.107167
R13103 VSS.n3130 VSS.n3129 0.107167
R13104 VSS.n3209 VSS.n3208 0.107167
R13105 VSS.n3288 VSS.n3287 0.107167
R13106 VSS.n2986 VSS.n2981 0.101624
R13107 VSS.n2990 VSS.n2986 0.101624
R13108 VSS.n2995 VSS.n2990 0.101624
R13109 VSS.n3000 VSS.n2995 0.101624
R13110 VSS.n3004 VSS.n3000 0.101624
R13111 VSS.n3009 VSS.n3004 0.101624
R13112 VSS.n3015 VSS.n3009 0.101624
R13113 VSS.n3020 VSS.n3015 0.101624
R13114 VSS.n3024 VSS.n3020 0.101624
R13115 VSS.n3029 VSS.n3024 0.101624
R13116 VSS.n3052 VSS.n3047 0.101624
R13117 VSS.n3056 VSS.n3052 0.101624
R13118 VSS.n3061 VSS.n3056 0.101624
R13119 VSS.n3065 VSS.n3061 0.101624
R13120 VSS.n3070 VSS.n3065 0.101624
R13121 VSS.n3074 VSS.n3070 0.101624
R13122 VSS.n3079 VSS.n3074 0.101624
R13123 VSS.n3103 VSS.n3099 0.101624
R13124 VSS.n3108 VSS.n3103 0.101624
R13125 VSS.n3112 VSS.n3108 0.101624
R13126 VSS.n3117 VSS.n3112 0.101624
R13127 VSS.n3121 VSS.n3117 0.101624
R13128 VSS.n3126 VSS.n3121 0.101624
R13129 VSS.n3131 VSS.n3126 0.101624
R13130 VSS.n3153 VSS.n3149 0.101624
R13131 VSS.n3158 VSS.n3153 0.101624
R13132 VSS.n3162 VSS.n3158 0.101624
R13133 VSS.n3167 VSS.n3162 0.101624
R13134 VSS.n3173 VSS.n3167 0.101624
R13135 VSS.n3178 VSS.n3173 0.101624
R13136 VSS.n3182 VSS.n3178 0.101624
R13137 VSS.n3205 VSS.n3200 0.101624
R13138 VSS.n3210 VSS.n3205 0.101624
R13139 VSS.n3214 VSS.n3210 0.101624
R13140 VSS.n3219 VSS.n3214 0.101624
R13141 VSS.n3223 VSS.n3219 0.101624
R13142 VSS.n3228 VSS.n3223 0.101624
R13143 VSS.n3232 VSS.n3228 0.101624
R13144 VSS.n3257 VSS.n3252 0.101624
R13145 VSS.n3261 VSS.n3257 0.101624
R13146 VSS.n3266 VSS.n3261 0.101624
R13147 VSS.n3270 VSS.n3266 0.101624
R13148 VSS.n3275 VSS.n3270 0.101624
R13149 VSS.n3279 VSS.n3275 0.101624
R13150 VSS.n3284 VSS.n3279 0.101624
R13151 VSS.n3307 VSS.n3302 0.101624
R13152 VSS.n3311 VSS.n3307 0.101624
R13153 VSS.n3316 VSS.n3311 0.101624
R13154 VSS.n3320 VSS.n3316 0.101624
R13155 VSS.n3325 VSS.n3320 0.101624
R13156 VSS.n3331 VSS.n3325 0.101624
R13157 VSS.n3336 VSS.n3331 0.101624
R13158 VSS.n3340 VSS.n3336 0.101624
R13159 VSS.n3345 VSS.n3340 0.101624
R13160 VSS.n3349 VSS.n3345 0.101624
R13161 VSS.n3354 VSS.n3349 0.101624
R13162 VSS.n3358 VSS.n3354 0.101624
R13163 VSS.n3365 VSS.n3358 0.101624
R13164 VSS.n3367 VSS.n3365 0.101624
R13165 VSS.n3369 VSS.n3367 0.101624
R13166 VSS.n3409 VSS.n3408 0.100111
R13167 VSS.n3404 VSS.n3403 0.100111
R13168 VSS.n551 VSS.n550 0.0974697
R13169 VSS.n730 VSS.n726 0.0974697
R13170 VSS.n740 VSS.n739 0.0974697
R13171 VSS.n754 VSS.n750 0.0974697
R13172 VSS.n261 VSS.n258 0.0971038
R13173 VSS.n412 VSS.n410 0.0971038
R13174 VSS.n432 VSS.n429 0.0971038
R13175 VSS.n475 VSS.n473 0.0971038
R13176 VSS.n489 VSS.n486 0.0971038
R13177 VSS.n501 VSS.n497 0.0971038
R13178 VSS.n846 VSS.n844 0.0971038
R13179 VSS.n860 VSS.n859 0.0971038
R13180 VSS.n863 VSS.n860 0.0971038
R13181 VSS.n969 VSS.n968 0.0971038
R13182 VSS.n1035 VSS.n1034 0.0971038
R13183 VSS.n1047 VSS.n1045 0.0971038
R13184 VSS.n1063 VSS.n1060 0.0971038
R13185 VSS.n1146 VSS.n1142 0.0971038
R13186 VSS.n1188 VSS.n1187 0.0971038
R13187 VSS.n1201 VSS.n1199 0.0971038
R13188 VSS.n1239 VSS.n1236 0.0971038
R13189 VSS.n1299 VSS.n1295 0.0971038
R13190 VSS.n1309 VSS.n1308 0.0971038
R13191 VSS.n1324 VSS.n1320 0.0971038
R13192 VSS.n1383 VSS.n1379 0.0971038
R13193 VSS.n1425 VSS.n1422 0.0971038
R13194 VSS.n1438 VSS.n1434 0.0971038
R13195 VSS.n1449 VSS.n1448 0.0971038
R13196 VSS.n1489 VSS.n1487 0.0971038
R13197 VSS.n1502 VSS.n1499 0.0971038
R13198 VSS.n1515 VSS.n1514 0.0971038
R13199 VSS.n1523 VSS.n1520 0.0971038
R13200 VSS.n1531 VSS.n1530 0.0971038
R13201 VSS.n1566 VSS.n1564 0.0971038
R13202 VSS.n1598 VSS.n1597 0.0971038
R13203 VSS.n3289 VSS.n3284 0.0964293
R13204 VSS.n2917 VSS.n2879 0.0959291
R13205 VSS.n3047 VSS.n3042 0.0860408
R13206 VSS.n3237 VSS.n3232 0.0860408
R13207 VSS.n2941 VSS.n2940 0.0855498
R13208 VSS.n204 VSS.n203 0.0833353
R13209 VSS.n191 VSS.n190 0.0830953
R13210 VSS.n375 VSS.n290 0.082675
R13211 VSS.n178 VSS.n177 0.0815709
R13212 VSS.n2930 VSS.n2926 0.0808571
R13213 VSS.n2934 VSS.n2930 0.0808571
R13214 VSS.n2938 VSS.n2934 0.0808571
R13215 VSS.n2945 VSS.n2938 0.0808571
R13216 VSS.n2949 VSS.n2945 0.0808571
R13217 VSS.n2953 VSS.n2949 0.0808571
R13218 VSS.n2957 VSS.n2953 0.0808571
R13219 VSS.n2961 VSS.n2957 0.0808571
R13220 VSS.n2965 VSS.n2961 0.0808571
R13221 VSS.n2969 VSS.n2965 0.0808571
R13222 VSS.n2973 VSS.n2969 0.0808571
R13223 VSS.n2975 VSS.n2973 0.0808571
R13224 VSS.n2976 VSS.n2975 0.0808571
R13225 VSS.n165 VSS.n164 0.0798057
R13226 VSS.n3099 VSS.n3094 0.0756524
R13227 VSS.n3187 VSS.n3182 0.0756524
R13228 VSS VSS.n3454 0.0715332
R13229 VSS.n2343 VSS.n2342 0.0700652
R13230 VSS.n2467 VSS.n2466 0.0700652
R13231 VSS.n2591 VSS.n2590 0.0700652
R13232 VSS.n2715 VSS.n2714 0.0700652
R13233 VSS.n2839 VSS.n2838 0.0700652
R13234 VSS.n3440 VSS.n3435 0.0692023
R13235 VSS.n3435 VSS.n3430 0.0692023
R13236 VSS.n3430 VSS.n3425 0.0692023
R13237 VSS.n3425 VSS.n3420 0.0692023
R13238 VSS.n3420 VSS.n3415 0.0692023
R13239 VSS.n3415 VSS.n3410 0.0692023
R13240 VSS.n3410 VSS.n3405 0.0692023
R13241 VSS.n3405 VSS.n3400 0.0692023
R13242 VSS.n3400 VSS.n3395 0.0692023
R13243 VSS.n3395 VSS.n3390 0.0692023
R13244 VSS.n3390 VSS.n3385 0.0692023
R13245 VSS.n3385 VSS.n3380 0.0692023
R13246 VSS.n3380 VSS.n3375 0.0692023
R13247 VSS.n3375 VSS.n3371 0.0692023
R13248 VSS.n3135 VSS.n3131 0.0652639
R13249 VSS.n3149 VSS.n3144 0.0652639
R13250 VSS.n1722 VSS.n1714 0.059284
R13251 VSS.n1731 VSS.n1723 0.059284
R13252 VSS.n1740 VSS.n1732 0.059284
R13253 VSS.n1749 VSS.n1741 0.059284
R13254 VSS.n1758 VSS.n1750 0.059284
R13255 VSS.n1767 VSS.n1759 0.059284
R13256 VSS.n1776 VSS.n1768 0.059284
R13257 VSS.n1785 VSS.n1777 0.059284
R13258 VSS.n1794 VSS.n1786 0.059284
R13259 VSS.n1803 VSS.n1795 0.059284
R13260 VSS.n1812 VSS.n1804 0.059284
R13261 VSS.n1821 VSS.n1813 0.059284
R13262 VSS.n1830 VSS.n1822 0.059284
R13263 VSS.n1839 VSS.n1831 0.059284
R13264 VSS.n1848 VSS.n1840 0.059284
R13265 VSS.n1857 VSS.n1849 0.059284
R13266 VSS.n1866 VSS.n1858 0.059284
R13267 VSS.n1875 VSS.n1867 0.059284
R13268 VSS.n1884 VSS.n1876 0.059284
R13269 VSS.n1901 VSS.n1893 0.059284
R13270 VSS.n1910 VSS.n1902 0.059284
R13271 VSS.n1919 VSS.n1911 0.059284
R13272 VSS.n1928 VSS.n1920 0.059284
R13273 VSS.n1937 VSS.n1929 0.059284
R13274 VSS.n1946 VSS.n1938 0.059284
R13275 VSS.n1955 VSS.n1947 0.059284
R13276 VSS.n1964 VSS.n1956 0.059284
R13277 VSS.n1973 VSS.n1965 0.059284
R13278 VSS.n1982 VSS.n1974 0.059284
R13279 VSS.n1991 VSS.n1983 0.059284
R13280 VSS.n2000 VSS.n1992 0.059284
R13281 VSS.n2009 VSS.n2001 0.059284
R13282 VSS.n2018 VSS.n2010 0.059284
R13283 VSS.n2027 VSS.n2019 0.059284
R13284 VSS.n2036 VSS.n2028 0.059284
R13285 VSS.n2045 VSS.n2037 0.059284
R13286 VSS.n2054 VSS.n2046 0.059284
R13287 VSS.n2063 VSS.n2055 0.059284
R13288 VSS.n2080 VSS.n2072 0.059284
R13289 VSS.n2089 VSS.n2081 0.059284
R13290 VSS.n2098 VSS.n2090 0.059284
R13291 VSS.n2107 VSS.n2099 0.059284
R13292 VSS.n2116 VSS.n2108 0.059284
R13293 VSS.n2125 VSS.n2117 0.059284
R13294 VSS.n2134 VSS.n2126 0.059284
R13295 VSS.n2143 VSS.n2135 0.059284
R13296 VSS.n2152 VSS.n2144 0.059284
R13297 VSS.n2161 VSS.n2153 0.059284
R13298 VSS.n2170 VSS.n2162 0.059284
R13299 VSS.n2179 VSS.n2171 0.059284
R13300 VSS.n2188 VSS.n2180 0.059284
R13301 VSS.n2197 VSS.n2189 0.059284
R13302 VSS.n2206 VSS.n2198 0.059284
R13303 VSS.n2215 VSS.n2207 0.059284
R13304 VSS.n2224 VSS.n2216 0.059284
R13305 VSS.n2233 VSS.n2225 0.059284
R13306 VSS.n2242 VSS.n2234 0.059284
R13307 VSS.n2286 VSS.n2276 0.0581923
R13308 VSS.n2292 VSS.n2286 0.0581923
R13309 VSS.n2300 VSS.n2292 0.0581923
R13310 VSS.n2306 VSS.n2300 0.0581923
R13311 VSS.n2314 VSS.n2306 0.0581923
R13312 VSS.n2320 VSS.n2314 0.0581923
R13313 VSS.n2330 VSS.n2320 0.0581923
R13314 VSS.n2336 VSS.n2330 0.0581923
R13315 VSS.n2344 VSS.n2336 0.0581923
R13316 VSS.n2351 VSS.n2344 0.0581923
R13317 VSS.n2358 VSS.n2351 0.0581923
R13318 VSS.n2365 VSS.n2358 0.0581923
R13319 VSS.n2372 VSS.n2365 0.0581923
R13320 VSS.n2379 VSS.n2372 0.0581923
R13321 VSS.n2386 VSS.n2379 0.0581923
R13322 VSS.n2424 VSS.n2416 0.0581923
R13323 VSS.n2430 VSS.n2424 0.0581923
R13324 VSS.n2438 VSS.n2430 0.0581923
R13325 VSS.n2444 VSS.n2438 0.0581923
R13326 VSS.n2454 VSS.n2444 0.0581923
R13327 VSS.n2460 VSS.n2454 0.0581923
R13328 VSS.n2468 VSS.n2460 0.0581923
R13329 VSS.n2475 VSS.n2468 0.0581923
R13330 VSS.n2503 VSS.n2496 0.0581923
R13331 VSS.n2510 VSS.n2503 0.0581923
R13332 VSS.n2518 VSS.n2510 0.0581923
R13333 VSS.n2524 VSS.n2518 0.0581923
R13334 VSS.n2534 VSS.n2524 0.0581923
R13335 VSS.n2540 VSS.n2534 0.0581923
R13336 VSS.n2548 VSS.n2540 0.0581923
R13337 VSS.n2554 VSS.n2548 0.0581923
R13338 VSS.n2584 VSS.n2578 0.0581923
R13339 VSS.n2592 VSS.n2584 0.0581923
R13340 VSS.n2599 VSS.n2592 0.0581923
R13341 VSS.n2606 VSS.n2599 0.0581923
R13342 VSS.n2613 VSS.n2606 0.0581923
R13343 VSS.n2620 VSS.n2613 0.0581923
R13344 VSS.n2627 VSS.n2620 0.0581923
R13345 VSS.n2634 VSS.n2627 0.0581923
R13346 VSS.n2672 VSS.n2664 0.0581923
R13347 VSS.n2678 VSS.n2672 0.0581923
R13348 VSS.n2686 VSS.n2678 0.0581923
R13349 VSS.n2692 VSS.n2686 0.0581923
R13350 VSS.n2702 VSS.n2692 0.0581923
R13351 VSS.n2708 VSS.n2702 0.0581923
R13352 VSS.n2716 VSS.n2708 0.0581923
R13353 VSS.n2751 VSS.n2744 0.0581923
R13354 VSS.n2758 VSS.n2751 0.0581923
R13355 VSS.n2766 VSS.n2758 0.0581923
R13356 VSS.n2772 VSS.n2766 0.0581923
R13357 VSS.n2782 VSS.n2772 0.0581923
R13358 VSS.n2788 VSS.n2782 0.0581923
R13359 VSS.n2796 VSS.n2788 0.0581923
R13360 VSS.n2832 VSS.n2826 0.0581923
R13361 VSS.n2840 VSS.n2832 0.0581923
R13362 VSS.n2847 VSS.n2840 0.0581923
R13363 VSS.n2854 VSS.n2847 0.0581923
R13364 VSS.n2861 VSS.n2854 0.0581923
R13365 VSS.n2868 VSS.n2861 0.0581923
R13366 VSS.n2875 VSS.n2868 0.0581923
R13367 VSS.n2879 VSS.n2875 0.0581923
R13368 VSS.n2394 VSS.n2386 0.056083
R13369 VSS.n107 VSS.n106 0.0549681
R13370 VSS.n106 VSS.n105 0.0549681
R13371 VSS.n3083 VSS.n3079 0.0548754
R13372 VSS.n3200 VSS.n3196 0.0548754
R13373 VSS.n2664 VSS.n2658 0.0546769
R13374 VSS.n2744 VSS.n2737 0.0490522
R13375 VSS.n562 VSS.n557 0.0489848
R13376 VSS.n562 VSS.n561 0.0489848
R13377 VSS.n576 VSS.n570 0.0489848
R13378 VSS.n585 VSS.n583 0.0489848
R13379 VSS.n696 VSS.n694 0.0489848
R13380 VSS.n763 VSS.n762 0.0489848
R13381 VSS.n333 VSS.n297 0.0488019
R13382 VSS.n227 VSS.n226 0.0488019
R13383 VSS.n1023 VSS.n1022 0.0488019
R13384 VSS.n1178 VSS.n1177 0.0488019
R13385 VSS.n1193 VSS.n1192 0.0488019
R13386 VSS.n1281 VSS.n1279 0.0488019
R13387 VSS.n1294 VSS.n1291 0.0488019
R13388 VSS.n1331 VSS.n1330 0.0488019
R13389 VSS.n1360 VSS.n1358 0.0488019
R13390 VSS.n1493 VSS.n1492 0.0488019
R13391 VSS.n1634 VSS.n1633 0.0488019
R13392 VSS.n3033 VSS.n3029 0.0444869
R13393 VSS.n3252 VSS.n3246 0.0444869
R13394 VSS.n2826 VSS.n2816 0.0434274
R13395 VSS.n647 VSS.n646 0.0361578
R13396 VSS.n382 VSS.n381 0.0345909
R13397 VSS.n385 VSS.n384 0.0345909
R13398 VSS.n399 VSS.n398 0.0345909
R13399 VSS.n402 VSS.n401 0.0345909
R13400 VSS.n446 VSS.n445 0.0345909
R13401 VSS.n449 VSS.n448 0.0345909
R13402 VSS.n464 VSS.n463 0.0345909
R13403 VSS.n467 VSS.n466 0.0345909
R13404 VSS.n600 VSS.n599 0.0345909
R13405 VSS.n604 VSS.n603 0.0345909
R13406 VSS.n618 VSS.n617 0.0345909
R13407 VSS.n622 VSS.n621 0.0345909
R13408 VSS.n631 VSS.n630 0.0345909
R13409 VSS.n634 VSS.n633 0.0345909
R13410 VSS.n650 VSS.n649 0.0345909
R13411 VSS.n918 VSS.n917 0.0345909
R13412 VSS.n921 VSS.n920 0.0345909
R13413 VSS.n935 VSS.n934 0.0345909
R13414 VSS.n938 VSS.n937 0.0345909
R13415 VSS.n1072 VSS.n1071 0.0345909
R13416 VSS.n1075 VSS.n1074 0.0345909
R13417 VSS.n1089 VSS.n1088 0.0345909
R13418 VSS.n1092 VSS.n1091 0.0345909
R13419 VSS.n1248 VSS.n1247 0.0345909
R13420 VSS.n1251 VSS.n1250 0.0345909
R13421 VSS.n1265 VSS.n1264 0.0345909
R13422 VSS.n1268 VSS.n1267 0.0345909
R13423 VSS.n1396 VSS.n1395 0.0345909
R13424 VSS.n1399 VSS.n1398 0.0345909
R13425 VSS.n1413 VSS.n1412 0.0345909
R13426 VSS.n1416 VSS.n1415 0.0345909
R13427 VSS.n1540 VSS.n1539 0.0345909
R13428 VSS.n1543 VSS.n1542 0.0345909
R13429 VSS.n1557 VSS.n1556 0.0345909
R13430 VSS.n1560 VSS.n1559 0.0345909
R13431 VSS.n1686 VSS.n1685 0.0345909
R13432 VSS.n1689 VSS.n1688 0.0345909
R13433 VSS.n3302 VSS.n3298 0.0340984
R13434 VSS.n2802 VSS.n2796 0.0335842
R13435 VSS.n207 VSS.n206 0.0292356
R13436 VSS.n2723 VSS.n2716 0.0279595
R13437 VSS.n1880 VSS.n1877 0.0278438
R13438 VSS.n1871 VSS.n1868 0.0278438
R13439 VSS.n1862 VSS.n1859 0.0278438
R13440 VSS.n1853 VSS.n1850 0.0278438
R13441 VSS.n1844 VSS.n1841 0.0278438
R13442 VSS.n1835 VSS.n1832 0.0278438
R13443 VSS.n1826 VSS.n1823 0.0278438
R13444 VSS.n1817 VSS.n1814 0.0278438
R13445 VSS.n1808 VSS.n1805 0.0278438
R13446 VSS.n1799 VSS.n1796 0.0278438
R13447 VSS.n1790 VSS.n1787 0.0278438
R13448 VSS.n1781 VSS.n1778 0.0278438
R13449 VSS.n1772 VSS.n1769 0.0278438
R13450 VSS.n1763 VSS.n1760 0.0278438
R13451 VSS.n1754 VSS.n1751 0.0278438
R13452 VSS.n1745 VSS.n1742 0.0278438
R13453 VSS.n1736 VSS.n1733 0.0278438
R13454 VSS.n1727 VSS.n1724 0.0278438
R13455 VSS.n1718 VSS.n1715 0.0278438
R13456 VSS.n1709 VSS.n1706 0.0278438
R13457 VSS.n2059 VSS.n2056 0.0278438
R13458 VSS.n2050 VSS.n2047 0.0278438
R13459 VSS.n2041 VSS.n2038 0.0278438
R13460 VSS.n2032 VSS.n2029 0.0278438
R13461 VSS.n2023 VSS.n2020 0.0278438
R13462 VSS.n2014 VSS.n2011 0.0278438
R13463 VSS.n2005 VSS.n2002 0.0278438
R13464 VSS.n1996 VSS.n1993 0.0278438
R13465 VSS.n1987 VSS.n1984 0.0278438
R13466 VSS.n1978 VSS.n1975 0.0278438
R13467 VSS.n1969 VSS.n1966 0.0278438
R13468 VSS.n1960 VSS.n1957 0.0278438
R13469 VSS.n1951 VSS.n1948 0.0278438
R13470 VSS.n1942 VSS.n1939 0.0278438
R13471 VSS.n1933 VSS.n1930 0.0278438
R13472 VSS.n1924 VSS.n1921 0.0278438
R13473 VSS.n1915 VSS.n1912 0.0278438
R13474 VSS.n1906 VSS.n1903 0.0278438
R13475 VSS.n1897 VSS.n1894 0.0278438
R13476 VSS.n1888 VSS.n1885 0.0278438
R13477 VSS.n2238 VSS.n2235 0.0278438
R13478 VSS.n2229 VSS.n2226 0.0278438
R13479 VSS.n2220 VSS.n2217 0.0278438
R13480 VSS.n2211 VSS.n2208 0.0278438
R13481 VSS.n2202 VSS.n2199 0.0278438
R13482 VSS.n2193 VSS.n2190 0.0278438
R13483 VSS.n2184 VSS.n2181 0.0278438
R13484 VSS.n2175 VSS.n2172 0.0278438
R13485 VSS.n2166 VSS.n2163 0.0278438
R13486 VSS.n2157 VSS.n2154 0.0278438
R13487 VSS.n2148 VSS.n2145 0.0278438
R13488 VSS.n2139 VSS.n2136 0.0278438
R13489 VSS.n2130 VSS.n2127 0.0278438
R13490 VSS.n2121 VSS.n2118 0.0278438
R13491 VSS.n2112 VSS.n2109 0.0278438
R13492 VSS.n2103 VSS.n2100 0.0278438
R13493 VSS.n2094 VSS.n2091 0.0278438
R13494 VSS.n2085 VSS.n2082 0.0278438
R13495 VSS.n2076 VSS.n2073 0.0278438
R13496 VSS.n2067 VSS.n2064 0.0278438
R13497 VSS.n194 VSS.n193 0.0277989
R13498 VSS.n181 VSS.n180 0.0277989
R13499 VSS.n154 VSS.n153 0.027734
R13500 VSS.n645 VSS.n644 0.0273716
R13501 VSS.n3445 VSS.n3440 0.0269538
R13502 VSS.n168 VSS.n167 0.0263621
R13503 VSS.n948 VSS.n947 0.0247248
R13504 VSS.n960 VSS.n959 0.0247248
R13505 VSS.n973 VSS.n972 0.0247248
R13506 VSS.n1006 VSS.n1005 0.0247248
R13507 VSS.n1016 VSS.n1015 0.0247248
R13508 VSS.n1027 VSS.n1026 0.0247248
R13509 VSS.n1040 VSS.n1039 0.0247248
R13510 VSS.n1104 VSS.n1103 0.0247248
R13511 VSS.n1139 VSS.n1138 0.0247248
R13512 VSS.n1150 VSS.n1149 0.0247248
R13513 VSS.n1160 VSS.n1159 0.0247248
R13514 VSS.n1171 VSS.n1170 0.0247248
R13515 VSS.n1182 VSS.n1181 0.0247248
R13516 VSS.n1197 VSS.n1196 0.0247248
R13517 VSS.n1277 VSS.n1276 0.0247248
R13518 VSS.n1289 VSS.n1288 0.0247248
R13519 VSS.n1303 VSS.n1302 0.0247248
R13520 VSS.n1313 VSS.n1312 0.0247248
R13521 VSS.n1327 VSS.n1326 0.0247248
R13522 VSS.n1335 VSS.n1334 0.0247248
R13523 VSS.n1367 VSS.n1366 0.0247248
R13524 VSS.n1429 VSS.n1428 0.0247248
R13525 VSS.n1442 VSS.n1441 0.0247248
R13526 VSS.n1454 VSS.n1453 0.0247248
R13527 VSS.n1464 VSS.n1463 0.0247248
R13528 VSS.n1485 VSS.n1484 0.0247248
R13529 VSS.n1497 VSS.n1496 0.0247248
R13530 VSS.n1510 VSS.n1509 0.0247248
R13531 VSS.n1571 VSS.n1570 0.0247248
R13532 VSS.n1581 VSS.n1580 0.0247248
R13533 VSS.n1602 VSS.n1601 0.0247248
R13534 VSS.n1613 VSS.n1612 0.0247248
R13535 VSS.n1628 VSS.n1627 0.0247248
R13536 VSS.n1638 VSS.n1637 0.0247248
R13537 VSS.n1651 VSS.n1650 0.0247248
R13538 VSS.n1674 VSS.n1673 0.0247248
R13539 VSS.n1669 VSS.n1668 0.0247248
R13540 VSS.n1701 VSS.n1700 0.0247248
R13541 VSS.n278 VSS.n277 0.0247248
R13542 VSS.n265 VSS.n264 0.0247248
R13543 VSS.n253 VSS.n252 0.0247248
R13544 VSS.n241 VSS.n240 0.0247248
R13545 VSS.n231 VSS.n230 0.0247248
R13546 VSS.n419 VSS.n418 0.0247248
R13547 VSS.n480 VSS.n479 0.0247248
R13548 VSS.n494 VSS.n493 0.0247248
R13549 VSS.n505 VSS.n504 0.0247248
R13550 VSS.n543 VSS.n542 0.0247248
R13551 VSS.n554 VSS.n553 0.0247248
R13552 VSS.n566 VSS.n565 0.0247248
R13553 VSS.n580 VSS.n579 0.0247248
R13554 VSS.n708 VSS.n707 0.0247248
R13555 VSS.n720 VSS.n719 0.0247248
R13556 VSS.n734 VSS.n733 0.0247248
R13557 VSS.n744 VSS.n743 0.0247248
R13558 VSS.n757 VSS.n756 0.0247248
R13559 VSS.n767 VSS.n766 0.0247248
R13560 VSS.n780 VSS.n779 0.0247248
R13561 VSS.n841 VSS.n840 0.0247248
R13562 VSS.n854 VSS.n853 0.0247248
R13563 VSS.n867 VSS.n866 0.0247248
R13564 VSS.n878 VSS.n877 0.0247248
R13565 VSS.n2919 VSS.n2917 0.0231131
R13566 VSS.n3449 VSS.n3445 0.0231131
R13567 VSS.n912 VSS.n911 0.0227868
R13568 VSS.n1066 VSS.n1065 0.0227868
R13569 VSS.n1242 VSS.n1241 0.0227868
R13570 VSS.n1390 VSS.n1389 0.0227868
R13571 VSS.n1534 VSS.n1533 0.0227868
R13572 VSS.n1680 VSS.n1679 0.0227868
R13573 VSS.n288 VSS.n287 0.0227868
R13574 VSS.n440 VSS.n439 0.0227868
R13575 VSS.n831 VSS.n828 0.0227868
R13576 VSS.n2642 VSS.n2634 0.0223348
R13577 VSS.n912 VSS.n903 0.0218178
R13578 VSS.n1066 VSS.n1057 0.0218178
R13579 VSS.n1242 VSS.n1208 0.0218178
R13580 VSS.n1390 VSS.n1384 0.0218178
R13581 VSS.n1534 VSS.n1525 0.0218178
R13582 VSS.n1680 VSS.n1663 0.0218178
R13583 VSS.n289 VSS.n288 0.0218178
R13584 VSS.n440 VSS.n434 0.0218178
R13585 VSS.n594 VSS.n593 0.0218178
R13586 VSS.n828 VSS.n827 0.0218178
R13587 VSS.n2416 VSS.n2410 0.0209286
R13588 VSS.n691 VSS.n657 0.0208704
R13589 VSS.n388 VSS.n387 0.0207922
R13590 VSS.n392 VSS.n391 0.0207922
R13591 VSS.n396 VSS.n395 0.0207922
R13592 VSS.n452 VSS.n451 0.0207922
R13593 VSS.n456 VSS.n455 0.0207922
R13594 VSS.n460 VSS.n459 0.0207922
R13595 VSS.n607 VSS.n606 0.0207922
R13596 VSS.n611 VSS.n610 0.0207922
R13597 VSS.n615 VSS.n614 0.0207922
R13598 VSS.n637 VSS.n636 0.0207922
R13599 VSS.n641 VSS.n640 0.0207922
R13600 VSS.n924 VSS.n923 0.0207922
R13601 VSS.n928 VSS.n927 0.0207922
R13602 VSS.n932 VSS.n931 0.0207922
R13603 VSS.n1078 VSS.n1077 0.0207922
R13604 VSS.n1082 VSS.n1081 0.0207922
R13605 VSS.n1086 VSS.n1085 0.0207922
R13606 VSS.n1254 VSS.n1253 0.0207922
R13607 VSS.n1258 VSS.n1257 0.0207922
R13608 VSS.n1262 VSS.n1261 0.0207922
R13609 VSS.n1402 VSS.n1401 0.0207922
R13610 VSS.n1406 VSS.n1405 0.0207922
R13611 VSS.n1410 VSS.n1409 0.0207922
R13612 VSS.n1546 VSS.n1545 0.0207922
R13613 VSS.n1550 VSS.n1549 0.0207922
R13614 VSS.n1554 VSS.n1553 0.0207922
R13615 VSS.n1692 VSS.n1691 0.0207922
R13616 VSS.n1699 VSS.n1698 0.0207922
R13617 VSS.n1005 VSS.n1004 0.0198798
R13618 VSS.n1015 VSS.n1014 0.0198798
R13619 VSS.n1159 VSS.n1158 0.0198798
R13620 VSS.n1170 VSS.n1169 0.0198798
R13621 VSS.n1312 VSS.n1311 0.0198798
R13622 VSS.n1326 VSS.n1325 0.0198798
R13623 VSS.n1463 VSS.n1462 0.0198798
R13624 VSS.n1484 VSS.n1483 0.0198798
R13625 VSS.n1612 VSS.n1611 0.0198798
R13626 VSS.n1627 VSS.n1626 0.0198798
R13627 VSS.n242 VSS.n241 0.0198798
R13628 VSS.n238 VSS.n231 0.0198798
R13629 VSS.n542 VSS.n541 0.0198798
R13630 VSS.n553 VSS.n552 0.0198798
R13631 VSS.n743 VSS.n742 0.0198798
R13632 VSS.n756 VSS.n755 0.0198798
R13633 VSS.n877 VSS.n876 0.0198798
R13634 VSS.n887 VSS.n886 0.0198798
R13635 VSS.n378 VSS.n377 0.0191688
R13636 VSS.n379 VSS.n378 0.0191688
R13637 VSS.n406 VSS.n405 0.0191688
R13638 VSS.n442 VSS.n441 0.0191688
R13639 VSS.n443 VSS.n442 0.0191688
R13640 VSS.n470 VSS.n469 0.0191688
R13641 VSS.n596 VSS.n595 0.0191688
R13642 VSS.n597 VSS.n596 0.0191688
R13643 VSS.n625 VSS.n624 0.0191688
R13644 VSS.n627 VSS.n626 0.0191688
R13645 VSS.n628 VSS.n627 0.0191688
R13646 VSS.n653 VSS.n652 0.0191688
R13647 VSS.n914 VSS.n913 0.0191688
R13648 VSS.n915 VSS.n914 0.0191688
R13649 VSS.n941 VSS.n940 0.0191688
R13650 VSS.n1068 VSS.n1067 0.0191688
R13651 VSS.n1069 VSS.n1068 0.0191688
R13652 VSS.n1095 VSS.n1094 0.0191688
R13653 VSS.n1244 VSS.n1243 0.0191688
R13654 VSS.n1245 VSS.n1244 0.0191688
R13655 VSS.n1271 VSS.n1270 0.0191688
R13656 VSS.n1392 VSS.n1391 0.0191688
R13657 VSS.n1393 VSS.n1392 0.0191688
R13658 VSS.n1419 VSS.n1418 0.0191688
R13659 VSS.n1536 VSS.n1535 0.0191688
R13660 VSS.n1537 VSS.n1536 0.0191688
R13661 VSS.n1563 VSS.n1562 0.0191688
R13662 VSS.n1682 VSS.n1681 0.0191688
R13663 VSS.n1683 VSS.n1682 0.0191688
R13664 VSS.n889 VSS.n888 0.0189109
R13665 VSS.n896 VSS.n890 0.0189109
R13666 VSS.n1003 VSS.n973 0.0189109
R13667 VSS.n1007 VSS.n1006 0.0189109
R13668 VSS.n1049 VSS.n1041 0.0189109
R13669 VSS.n1157 VSS.n1150 0.0189109
R13670 VSS.n1161 VSS.n1160 0.0189109
R13671 VSS.n1203 VSS.n1198 0.0189109
R13672 VSS.n1310 VSS.n1303 0.0189109
R13673 VSS.n1314 VSS.n1313 0.0189109
R13674 VSS.n1373 VSS.n1368 0.0189109
R13675 VSS.n1461 VSS.n1454 0.0189109
R13676 VSS.n1465 VSS.n1464 0.0189109
R13677 VSS.n1517 VSS.n1511 0.0189109
R13678 VSS.n1610 VSS.n1602 0.0189109
R13679 VSS.n1614 VSS.n1613 0.0189109
R13680 VSS.n1658 VSS.n1652 0.0189109
R13681 VSS.n1695 VSS.n1694 0.0189109
R13682 VSS.n1703 VSS.n1701 0.0189109
R13683 VSS.n252 VSS.n251 0.0189109
R13684 VSS.n240 VSS.n239 0.0189109
R13685 VSS.n423 VSS.n420 0.0189109
R13686 VSS.n540 VSS.n505 0.0189109
R13687 VSS.n544 VSS.n543 0.0189109
R13688 VSS.n586 VSS.n581 0.0189109
R13689 VSS.n741 VSS.n734 0.0189109
R13690 VSS.n745 VSS.n744 0.0189109
R13691 VSS.n787 VSS.n781 0.0189109
R13692 VSS.n875 VSS.n867 0.0189109
R13693 VSS.n879 VSS.n878 0.0189109
R13694 VSS.n199 VSS.n198 0.0187927
R13695 VSS.n648 VSS.n647 0.0185586
R13696 VSS.n377 VSS.n376 0.0183571
R13697 VSS.n441 VSS.n406 0.0183571
R13698 VSS.n595 VSS.n470 0.0183571
R13699 VSS.n626 VSS.n625 0.0183571
R13700 VSS.n913 VSS.n653 0.0183571
R13701 VSS.n1067 VSS.n941 0.0183571
R13702 VSS.n1243 VSS.n1095 0.0183571
R13703 VSS.n1391 VSS.n1271 0.0183571
R13704 VSS.n1535 VSS.n1419 0.0183571
R13705 VSS.n1681 VSS.n1563 0.0183571
R13706 VSS.n946 VSS.n945 0.0179419
R13707 VSS.n1275 VSS.n1274 0.0179419
R13708 VSS.n1427 VSS.n1426 0.0179419
R13709 VSS.n1569 VSS.n1568 0.0179419
R13710 VSS.n1676 VSS.n1675 0.0179419
R13711 VSS.n284 VSS.n279 0.0179419
R13712 VSS.n478 VSS.n477 0.0179419
R13713 VSS.n706 VSS.n705 0.0179419
R13714 VSS.n839 VSS.n838 0.0179419
R13715 VSS.n186 VSS.n185 0.0172683
R13716 VSS.n391 VSS.n390 0.0167338
R13717 VSS.n395 VSS.n394 0.0167338
R13718 VSS.n455 VSS.n454 0.0167338
R13719 VSS.n459 VSS.n458 0.0167338
R13720 VSS.n610 VSS.n609 0.0167338
R13721 VSS.n614 VSS.n613 0.0167338
R13722 VSS.n640 VSS.n639 0.0167338
R13723 VSS.n644 VSS.n643 0.0167338
R13724 VSS.n927 VSS.n926 0.0167338
R13725 VSS.n931 VSS.n930 0.0167338
R13726 VSS.n1081 VSS.n1080 0.0167338
R13727 VSS.n1085 VSS.n1084 0.0167338
R13728 VSS.n1257 VSS.n1256 0.0167338
R13729 VSS.n1261 VSS.n1260 0.0167338
R13730 VSS.n1405 VSS.n1404 0.0167338
R13731 VSS.n1409 VSS.n1408 0.0167338
R13732 VSS.n1549 VSS.n1548 0.0167338
R13733 VSS.n1553 VSS.n1552 0.0167338
R13734 VSS.n1698 VSS.n1697 0.0167338
R13735 VSS.n2562 VSS.n2554 0.0167101
R13736 VSS.n888 VSS.n655 0.0162407
R13737 VSS.n972 VSS.n971 0.0160039
R13738 VSS.n1026 VSS.n1025 0.0160039
R13739 VSS.n1149 VSS.n1148 0.0160039
R13740 VSS.n1181 VSS.n1180 0.0160039
R13741 VSS.n1302 VSS.n1301 0.0160039
R13742 VSS.n1334 VSS.n1333 0.0160039
R13743 VSS.n1496 VSS.n1495 0.0160039
R13744 VSS.n1601 VSS.n1600 0.0160039
R13745 VSS.n1637 VSS.n1636 0.0160039
R13746 VSS.n1665 VSS.n1664 0.0160039
R13747 VSS.n254 VSS.n253 0.0160039
R13748 VSS.n209 VSS.n208 0.0160039
R13749 VSS.n504 VSS.n503 0.0160039
R13750 VSS.n565 VSS.n564 0.0160039
R13751 VSS.n733 VSS.n732 0.0160039
R13752 VSS.n766 VSS.n765 0.0160039
R13753 VSS.n866 VSS.n865 0.0160039
R13754 VSS.n389 VSS.n388 0.0159221
R13755 VSS.n393 VSS.n392 0.0159221
R13756 VSS.n453 VSS.n452 0.0159221
R13757 VSS.n457 VSS.n456 0.0159221
R13758 VSS.n469 VSS.n468 0.0159221
R13759 VSS.n608 VSS.n607 0.0159221
R13760 VSS.n612 VSS.n611 0.0159221
R13761 VSS.n624 VSS.n623 0.0159221
R13762 VSS.n638 VSS.n637 0.0159221
R13763 VSS.n642 VSS.n641 0.0159221
R13764 VSS.n652 VSS.n651 0.0159221
R13765 VSS.n925 VSS.n924 0.0159221
R13766 VSS.n929 VSS.n928 0.0159221
R13767 VSS.n940 VSS.n939 0.0159221
R13768 VSS.n1079 VSS.n1078 0.0159221
R13769 VSS.n1083 VSS.n1082 0.0159221
R13770 VSS.n1094 VSS.n1093 0.0159221
R13771 VSS.n1255 VSS.n1254 0.0159221
R13772 VSS.n1259 VSS.n1258 0.0159221
R13773 VSS.n1270 VSS.n1269 0.0159221
R13774 VSS.n1403 VSS.n1402 0.0159221
R13775 VSS.n1407 VSS.n1406 0.0159221
R13776 VSS.n1418 VSS.n1417 0.0159221
R13777 VSS.n1547 VSS.n1546 0.0159221
R13778 VSS.n1551 VSS.n1550 0.0159221
R13779 VSS.n1562 VSS.n1561 0.0159221
R13780 VSS.n1693 VSS.n1692 0.0159221
R13781 VSS.n1704 VSS.n1699 0.0159221
R13782 VSS.n3450 VSS.n3449 0.0158894
R13783 VSS.n173 VSS.n172 0.0157439
R13784 VSS.n2496 VSS.n2489 0.0153039
R13785 VSS.n380 VSS.n379 0.0151104
R13786 VSS.n444 VSS.n443 0.0151104
R13787 VSS.n598 VSS.n597 0.0151104
R13788 VSS.n629 VSS.n628 0.0151104
R13789 VSS.n916 VSS.n915 0.0151104
R13790 VSS.n1070 VSS.n1069 0.0151104
R13791 VSS.n1246 VSS.n1245 0.0151104
R13792 VSS.n1394 VSS.n1393 0.0151104
R13793 VSS.n1538 VSS.n1537 0.0151104
R13794 VSS.n1684 VSS.n1683 0.0151104
R13795 VSS.n961 VSS.n960 0.0150349
R13796 VSS.n1017 VSS.n1016 0.0150349
R13797 VSS.n1037 VSS.n1028 0.0150349
R13798 VSS.n1140 VSS.n1139 0.0150349
R13799 VSS.n1172 VSS.n1171 0.0150349
R13800 VSS.n1194 VSS.n1183 0.0150349
R13801 VSS.n1290 VSS.n1289 0.0150349
R13802 VSS.n1328 VSS.n1327 0.0150349
R13803 VSS.n1364 VSS.n1336 0.0150349
R13804 VSS.n1443 VSS.n1442 0.0150349
R13805 VSS.n1486 VSS.n1485 0.0150349
R13806 VSS.n1507 VSS.n1498 0.0150349
R13807 VSS.n1582 VSS.n1581 0.0150349
R13808 VSS.n1629 VSS.n1628 0.0150349
R13809 VSS.n1648 VSS.n1639 0.0150349
R13810 VSS.n1668 VSS.n1667 0.0150349
R13811 VSS.n264 VSS.n263 0.0150349
R13812 VSS.n230 VSS.n229 0.0150349
R13813 VSS.n416 VSS.n408 0.0150349
R13814 VSS.n495 VSS.n494 0.0150349
R13815 VSS.n555 VSS.n554 0.0150349
R13816 VSS.n577 VSS.n567 0.0150349
R13817 VSS.n721 VSS.n720 0.0150349
R13818 VSS.n758 VSS.n757 0.0150349
R13819 VSS.n777 VSS.n768 0.0150349
R13820 VSS.n855 VSS.n854 0.0150349
R13821 VSS.n958 VSS.n957 0.0140659
R13822 VSS.n1137 VSS.n1136 0.0140659
R13823 VSS.n1287 VSS.n1286 0.0140659
R13824 VSS.n1440 VSS.n1439 0.0140659
R13825 VSS.n1579 VSS.n1578 0.0140659
R13826 VSS.n1671 VSS.n1670 0.0140659
R13827 VSS.n275 VSS.n266 0.0140659
R13828 VSS.n492 VSS.n491 0.0140659
R13829 VSS.n718 VSS.n717 0.0140659
R13830 VSS.n852 VSS.n851 0.0140659
R13831 VSS.n387 VSS.n386 0.013487
R13832 VSS.n451 VSS.n450 0.013487
R13833 VSS.n606 VSS.n605 0.013487
R13834 VSS.n636 VSS.n635 0.013487
R13835 VSS.n923 VSS.n922 0.013487
R13836 VSS.n1077 VSS.n1076 0.013487
R13837 VSS.n1253 VSS.n1252 0.013487
R13838 VSS.n1401 VSS.n1400 0.013487
R13839 VSS.n1545 VSS.n1544 0.013487
R13840 VSS.n1691 VSS.n1690 0.013487
R13841 VSS.n163 VSS.n160 0.0126951
R13842 VSS.n160 VSS.n159 0.0126951
R13843 VSS.n397 VSS.n396 0.0126753
R13844 VSS.n401 VSS.n400 0.0126753
R13845 VSS.n466 VSS.n465 0.0126753
R13846 VSS.n616 VSS.n615 0.0126753
R13847 VSS.n621 VSS.n620 0.0126753
R13848 VSS.n649 VSS.n648 0.0126753
R13849 VSS.n933 VSS.n932 0.0126753
R13850 VSS.n937 VSS.n936 0.0126753
R13851 VSS.n1087 VSS.n1086 0.0126753
R13852 VSS.n1091 VSS.n1090 0.0126753
R13853 VSS.n1263 VSS.n1262 0.0126753
R13854 VSS.n1267 VSS.n1266 0.0126753
R13855 VSS.n1411 VSS.n1410 0.0126753
R13856 VSS.n1415 VSS.n1414 0.0126753
R13857 VSS.n1555 VSS.n1554 0.0126753
R13858 VSS.n1559 VSS.n1558 0.0126753
R13859 VSS.n1705 VSS.n1704 0.0123316
R13860 VSS.n959 VSS.n958 0.0121279
R13861 VSS.n1039 VSS.n1038 0.0121279
R13862 VSS.n1138 VSS.n1137 0.0121279
R13863 VSS.n1196 VSS.n1195 0.0121279
R13864 VSS.n1288 VSS.n1287 0.0121279
R13865 VSS.n1366 VSS.n1365 0.0121279
R13866 VSS.n1441 VSS.n1440 0.0121279
R13867 VSS.n1509 VSS.n1508 0.0121279
R13868 VSS.n1580 VSS.n1579 0.0121279
R13869 VSS.n1650 VSS.n1649 0.0121279
R13870 VSS.n1670 VSS.n1669 0.0121279
R13871 VSS.n266 VSS.n265 0.0121279
R13872 VSS.n418 VSS.n417 0.0121279
R13873 VSS.n493 VSS.n492 0.0121279
R13874 VSS.n579 VSS.n578 0.0121279
R13875 VSS.n719 VSS.n718 0.0121279
R13876 VSS.n779 VSS.n778 0.0121279
R13877 VSS.n853 VSS.n852 0.0121279
R13878 VSS.n167 VSS.n166 0.0119943
R13879 VSS.n383 VSS.n382 0.0118636
R13880 VSS.n447 VSS.n446 0.0118636
R13881 VSS.n632 VSS.n631 0.0118636
R13882 VSS.n919 VSS.n918 0.0118636
R13883 VSS.n1073 VSS.n1072 0.0118636
R13884 VSS.n1249 VSS.n1248 0.0118636
R13885 VSS.n1397 VSS.n1396 0.0118636
R13886 VSS.n1541 VSS.n1540 0.0118636
R13887 VSS.n1687 VSS.n1686 0.0118636
R13888 VSS.n949 VSS.n948 0.0111589
R13889 VSS.n1024 VSS.n1017 0.0111589
R13890 VSS.n1028 VSS.n1027 0.0111589
R13891 VSS.n1105 VSS.n1104 0.0111589
R13892 VSS.n1179 VSS.n1172 0.0111589
R13893 VSS.n1183 VSS.n1182 0.0111589
R13894 VSS.n1278 VSS.n1277 0.0111589
R13895 VSS.n1332 VSS.n1328 0.0111589
R13896 VSS.n1336 VSS.n1335 0.0111589
R13897 VSS.n1430 VSS.n1429 0.0111589
R13898 VSS.n1494 VSS.n1486 0.0111589
R13899 VSS.n1498 VSS.n1497 0.0111589
R13900 VSS.n1572 VSS.n1571 0.0111589
R13901 VSS.n1635 VSS.n1629 0.0111589
R13902 VSS.n1639 VSS.n1638 0.0111589
R13903 VSS.n1673 VSS.n1672 0.0111589
R13904 VSS.n277 VSS.n276 0.0111589
R13905 VSS.n229 VSS.n228 0.0111589
R13906 VSS.n408 VSS.n407 0.0111589
R13907 VSS.n481 VSS.n480 0.0111589
R13908 VSS.n563 VSS.n555 0.0111589
R13909 VSS.n567 VSS.n566 0.0111589
R13910 VSS.n709 VSS.n708 0.0111589
R13911 VSS.n764 VSS.n758 0.0111589
R13912 VSS.n768 VSS.n767 0.0111589
R13913 VSS.n842 VSS.n841 0.0111589
R13914 VSS.n2482 VSS.n2475 0.0110854
R13915 VSS.n405 VSS.n404 0.0110519
R13916 VSS.n384 VSS.n383 0.0102403
R13917 VSS.n448 VSS.n447 0.0102403
R13918 VSS.n603 VSS.n602 0.0102403
R13919 VSS.n633 VSS.n632 0.0102403
R13920 VSS.n920 VSS.n919 0.0102403
R13921 VSS.n1074 VSS.n1073 0.0102403
R13922 VSS.n1250 VSS.n1249 0.0102403
R13923 VSS.n1398 VSS.n1397 0.0102403
R13924 VSS.n1542 VSS.n1541 0.0102403
R13925 VSS.n1688 VSS.n1687 0.0102403
R13926 VSS.n903 VSS.n898 0.0101899
R13927 VSS.n971 VSS.n970 0.0101899
R13928 VSS.n1057 VSS.n1051 0.0101899
R13929 VSS.n1102 VSS.n1101 0.0101899
R13930 VSS.n1148 VSS.n1147 0.0101899
R13931 VSS.n1208 VSS.n1205 0.0101899
R13932 VSS.n1301 VSS.n1300 0.0101899
R13933 VSS.n1384 VSS.n1375 0.0101899
R13934 VSS.n1451 VSS.n1450 0.0101899
R13935 VSS.n1525 VSS.n1519 0.0101899
R13936 VSS.n1600 VSS.n1599 0.0101899
R13937 VSS.n1663 VSS.n1660 0.0101899
R13938 VSS.n1677 VSS.n1676 0.0101899
R13939 VSS.n1666 VSS.n1665 0.0101899
R13940 VSS.n290 VSS.n289 0.0101899
R13941 VSS.n285 VSS.n284 0.0101899
R13942 VSS.n262 VSS.n254 0.0101899
R13943 VSS.n434 VSS.n425 0.0101899
R13944 VSS.n503 VSS.n502 0.0101899
R13945 VSS.n593 VSS.n588 0.0101899
R13946 VSS.n705 VSS.n699 0.0101899
R13947 VSS.n732 VSS.n731 0.0101899
R13948 VSS.n827 VSS.n789 0.0101899
R13949 VSS.n838 VSS.n833 0.0101899
R13950 VSS.n865 VSS.n864 0.0101899
R13951 VSS.n2578 VSS.n2568 0.00967918
R13952 VSS.n176 VSS.n173 0.00964634
R13953 VSS.n398 VSS.n397 0.00942857
R13954 VSS.n400 VSS.n399 0.00942857
R13955 VSS.n463 VSS.n462 0.00942857
R13956 VSS.n465 VSS.n464 0.00942857
R13957 VSS.n617 VSS.n616 0.00942857
R13958 VSS.n934 VSS.n933 0.00942857
R13959 VSS.n936 VSS.n935 0.00942857
R13960 VSS.n1088 VSS.n1087 0.00942857
R13961 VSS.n1090 VSS.n1089 0.00942857
R13962 VSS.n1264 VSS.n1263 0.00942857
R13963 VSS.n1266 VSS.n1265 0.00942857
R13964 VSS.n1412 VSS.n1411 0.00942857
R13965 VSS.n1414 VSS.n1413 0.00942857
R13966 VSS.n1556 VSS.n1555 0.00942857
R13967 VSS.n1558 VSS.n1557 0.00942857
R13968 VSS.n897 VSS.n896 0.00922093
R13969 VSS.n911 VSS.n905 0.00922093
R13970 VSS.n1050 VSS.n1049 0.00922093
R13971 VSS.n1065 VSS.n1059 0.00922093
R13972 VSS.n1204 VSS.n1203 0.00922093
R13973 VSS.n1241 VSS.n1210 0.00922093
R13974 VSS.n1374 VSS.n1373 0.00922093
R13975 VSS.n1389 VSS.n1386 0.00922093
R13976 VSS.n1452 VSS.n1451 0.00922093
R13977 VSS.n1518 VSS.n1517 0.00922093
R13978 VSS.n1533 VSS.n1527 0.00922093
R13979 VSS.n1659 VSS.n1658 0.00922093
R13980 VSS.n1679 VSS.n1678 0.00922093
R13981 VSS.n287 VSS.n286 0.00922093
R13982 VSS.n424 VSS.n423 0.00922093
R13983 VSS.n439 VSS.n436 0.00922093
R13984 VSS.n587 VSS.n586 0.00922093
R13985 VSS.n698 VSS.n697 0.00922093
R13986 VSS.n788 VSS.n787 0.00922093
R13987 VSS.n832 VSS.n831 0.00922093
R13988 VSS.n180 VSS.n179 0.00912069
R13989 VSS.n386 VSS.n385 0.00861688
R13990 VSS.n450 VSS.n449 0.00861688
R13991 VSS.n602 VSS.n601 0.00861688
R13992 VSS.n605 VSS.n604 0.00861688
R13993 VSS.n635 VSS.n634 0.00861688
R13994 VSS.n922 VSS.n921 0.00861688
R13995 VSS.n1076 VSS.n1075 0.00861688
R13996 VSS.n1252 VSS.n1251 0.00861688
R13997 VSS.n1400 VSS.n1399 0.00861688
R13998 VSS.n1544 VSS.n1543 0.00861688
R13999 VSS.n1690 VSS.n1689 0.00861688
R14000 VSS.n947 VSS.n946 0.00825194
R14001 VSS.n1101 VSS.n1100 0.00825194
R14002 VSS.n1103 VSS.n1102 0.00825194
R14003 VSS.n1276 VSS.n1275 0.00825194
R14004 VSS.n1428 VSS.n1427 0.00825194
R14005 VSS.n1570 VSS.n1569 0.00825194
R14006 VSS.n1675 VSS.n1674 0.00825194
R14007 VSS.n279 VSS.n278 0.00825194
R14008 VSS.n479 VSS.n478 0.00825194
R14009 VSS.n707 VSS.n706 0.00825194
R14010 VSS.n840 VSS.n839 0.00825194
R14011 VSS.n3038 VSS.n3033 0.00812712
R14012 VSS.n3042 VSS.n3038 0.00812712
R14013 VSS.n3088 VSS.n3083 0.00812712
R14014 VSS.n3094 VSS.n3088 0.00812712
R14015 VSS.n3140 VSS.n3135 0.00812712
R14016 VSS.n3144 VSS.n3140 0.00812712
R14017 VSS.n3191 VSS.n3187 0.00812712
R14018 VSS.n3196 VSS.n3191 0.00812712
R14019 VSS.n3241 VSS.n3237 0.00812712
R14020 VSS.n3246 VSS.n3241 0.00812712
R14021 VSS.n3293 VSS.n3289 0.00812712
R14022 VSS.n3298 VSS.n3293 0.00812712
R14023 VSS.n189 VSS.n186 0.00812195
R14024 VSS.n462 VSS.n461 0.00780519
R14025 VSS.n620 VSS.n619 0.00780519
R14026 VSS.n3450 VSS.n2919 0.00772362
R14027 VSS.n193 VSS.n192 0.00768391
R14028 VSS.n2400 VSS.n2394 0.00756991
R14029 VSS.n2410 VSS.n2400 0.00756991
R14030 VSS.n2489 VSS.n2482 0.00756991
R14031 VSS.n2568 VSS.n2562 0.00756991
R14032 VSS.n2648 VSS.n2642 0.00756991
R14033 VSS.n2658 VSS.n2648 0.00756991
R14034 VSS.n2730 VSS.n2723 0.00756991
R14035 VSS.n2737 VSS.n2730 0.00756991
R14036 VSS.n2810 VSS.n2802 0.00756991
R14037 VSS.n2816 VSS.n2810 0.00756991
R14038 VSS.n890 VSS.n889 0.00728295
R14039 VSS.n1041 VSS.n1040 0.00728295
R14040 VSS.n1198 VSS.n1197 0.00728295
R14041 VSS.n1368 VSS.n1367 0.00728295
R14042 VSS.n1453 VSS.n1452 0.00728295
R14043 VSS.n1511 VSS.n1510 0.00728295
R14044 VSS.n1652 VSS.n1651 0.00728295
R14045 VSS.n420 VSS.n419 0.00728295
R14046 VSS.n581 VSS.n580 0.00728295
R14047 VSS.n781 VSS.n780 0.00728295
R14048 VSS.n888 VSS.n887 0.00728295
R14049 VSS.n646 VSS.n645 0.00707944
R14050 VSS.n381 VSS.n380 0.00699351
R14051 VSS.n445 VSS.n444 0.00699351
R14052 VSS.n599 VSS.n598 0.00699351
R14053 VSS.n630 VSS.n629 0.00699351
R14054 VSS.n917 VSS.n916 0.00699351
R14055 VSS.n1071 VSS.n1070 0.00699351
R14056 VSS.n1247 VSS.n1246 0.00699351
R14057 VSS.n1395 VSS.n1394 0.00699351
R14058 VSS.n1539 VSS.n1538 0.00699351
R14059 VSS.n1685 VSS.n1684 0.00699351
R14060 VSS.n202 VSS.n199 0.00659756
R14061 VSS.n1883 VSS.n1880 0.00635938
R14062 VSS.n1874 VSS.n1871 0.00635938
R14063 VSS.n1865 VSS.n1862 0.00635938
R14064 VSS.n1856 VSS.n1853 0.00635938
R14065 VSS.n1847 VSS.n1844 0.00635938
R14066 VSS.n1838 VSS.n1835 0.00635938
R14067 VSS.n1829 VSS.n1826 0.00635938
R14068 VSS.n1820 VSS.n1817 0.00635938
R14069 VSS.n1811 VSS.n1808 0.00635938
R14070 VSS.n1802 VSS.n1799 0.00635938
R14071 VSS.n1793 VSS.n1790 0.00635938
R14072 VSS.n1784 VSS.n1781 0.00635938
R14073 VSS.n1775 VSS.n1772 0.00635938
R14074 VSS.n1766 VSS.n1763 0.00635938
R14075 VSS.n1757 VSS.n1754 0.00635938
R14076 VSS.n1748 VSS.n1745 0.00635938
R14077 VSS.n1739 VSS.n1736 0.00635938
R14078 VSS.n1730 VSS.n1727 0.00635938
R14079 VSS.n1721 VSS.n1718 0.00635938
R14080 VSS.n1712 VSS.n1709 0.00635938
R14081 VSS.n2062 VSS.n2059 0.00635938
R14082 VSS.n2053 VSS.n2050 0.00635938
R14083 VSS.n2044 VSS.n2041 0.00635938
R14084 VSS.n2035 VSS.n2032 0.00635938
R14085 VSS.n2026 VSS.n2023 0.00635938
R14086 VSS.n2017 VSS.n2014 0.00635938
R14087 VSS.n2008 VSS.n2005 0.00635938
R14088 VSS.n1999 VSS.n1996 0.00635938
R14089 VSS.n1990 VSS.n1987 0.00635938
R14090 VSS.n1981 VSS.n1978 0.00635938
R14091 VSS.n1972 VSS.n1969 0.00635938
R14092 VSS.n1963 VSS.n1960 0.00635938
R14093 VSS.n1954 VSS.n1951 0.00635938
R14094 VSS.n1945 VSS.n1942 0.00635938
R14095 VSS.n1936 VSS.n1933 0.00635938
R14096 VSS.n1927 VSS.n1924 0.00635938
R14097 VSS.n1918 VSS.n1915 0.00635938
R14098 VSS.n1909 VSS.n1906 0.00635938
R14099 VSS.n1900 VSS.n1897 0.00635938
R14100 VSS.n1891 VSS.n1888 0.00635938
R14101 VSS.n2241 VSS.n2238 0.00635938
R14102 VSS.n2232 VSS.n2229 0.00635938
R14103 VSS.n2223 VSS.n2220 0.00635938
R14104 VSS.n2214 VSS.n2211 0.00635938
R14105 VSS.n2205 VSS.n2202 0.00635938
R14106 VSS.n2196 VSS.n2193 0.00635938
R14107 VSS.n2187 VSS.n2184 0.00635938
R14108 VSS.n2178 VSS.n2175 0.00635938
R14109 VSS.n2169 VSS.n2166 0.00635938
R14110 VSS.n2160 VSS.n2157 0.00635938
R14111 VSS.n2151 VSS.n2148 0.00635938
R14112 VSS.n2142 VSS.n2139 0.00635938
R14113 VSS.n2133 VSS.n2130 0.00635938
R14114 VSS.n2124 VSS.n2121 0.00635938
R14115 VSS.n2115 VSS.n2112 0.00635938
R14116 VSS.n2106 VSS.n2103 0.00635938
R14117 VSS.n2097 VSS.n2094 0.00635938
R14118 VSS.n2088 VSS.n2085 0.00635938
R14119 VSS.n2079 VSS.n2076 0.00635938
R14120 VSS.n2070 VSS.n2067 0.00635938
R14121 VSS.n957 VSS.n949 0.00631395
R14122 VSS.n1136 VSS.n1105 0.00631395
R14123 VSS.n1286 VSS.n1278 0.00631395
R14124 VSS.n1439 VSS.n1430 0.00631395
R14125 VSS.n1578 VSS.n1572 0.00631395
R14126 VSS.n1672 VSS.n1671 0.00631395
R14127 VSS.n276 VSS.n275 0.00631395
R14128 VSS.n491 VSS.n481 0.00631395
R14129 VSS.n717 VSS.n709 0.00631395
R14130 VSS.n851 VSS.n842 0.00631395
R14131 VSS.n206 VSS.n205 0.00624713
R14132 VSS.n403 VSS.n402 0.00618182
R14133 VSS.n468 VSS.n467 0.00618182
R14134 VSS.n623 VSS.n622 0.00618182
R14135 VSS.n651 VSS.n650 0.00618182
R14136 VSS.n939 VSS.n938 0.00618182
R14137 VSS.n1093 VSS.n1092 0.00618182
R14138 VSS.n1269 VSS.n1268 0.00618182
R14139 VSS.n1417 VSS.n1416 0.00618182
R14140 VSS.n1561 VSS.n1560 0.00618182
R14141 VSS.n404 VSS.n403 0.00537013
R14142 VSS.n461 VSS.n460 0.00537013
R14143 VSS.n1038 VSS.n1037 0.00534496
R14144 VSS.n1195 VSS.n1194 0.00534496
R14145 VSS.n1365 VSS.n1364 0.00534496
R14146 VSS.n1508 VSS.n1507 0.00534496
R14147 VSS.n1649 VSS.n1648 0.00534496
R14148 VSS.n417 VSS.n416 0.00534496
R14149 VSS.n578 VSS.n577 0.00534496
R14150 VSS.n778 VSS.n777 0.00534496
R14151 VSS.n898 VSS.n897 0.00437597
R14152 VSS.n905 VSS.n904 0.00437597
R14153 VSS.n1004 VSS.n1003 0.00437597
R14154 VSS.n1014 VSS.n1007 0.00437597
R14155 VSS.n1051 VSS.n1050 0.00437597
R14156 VSS.n1059 VSS.n1058 0.00437597
R14157 VSS.n1158 VSS.n1157 0.00437597
R14158 VSS.n1169 VSS.n1161 0.00437597
R14159 VSS.n1205 VSS.n1204 0.00437597
R14160 VSS.n1210 VSS.n1209 0.00437597
R14161 VSS.n1311 VSS.n1310 0.00437597
R14162 VSS.n1325 VSS.n1314 0.00437597
R14163 VSS.n1375 VSS.n1374 0.00437597
R14164 VSS.n1386 VSS.n1385 0.00437597
R14165 VSS.n1462 VSS.n1461 0.00437597
R14166 VSS.n1483 VSS.n1465 0.00437597
R14167 VSS.n1519 VSS.n1518 0.00437597
R14168 VSS.n1527 VSS.n1526 0.00437597
R14169 VSS.n1611 VSS.n1610 0.00437597
R14170 VSS.n1626 VSS.n1614 0.00437597
R14171 VSS.n1660 VSS.n1659 0.00437597
R14172 VSS.n1678 VSS.n1677 0.00437597
R14173 VSS.n1696 VSS.n1695 0.00437597
R14174 VSS.n1703 VSS.n1702 0.00437597
R14175 VSS.n286 VSS.n285 0.00437597
R14176 VSS.n251 VSS.n242 0.00437597
R14177 VSS.n239 VSS.n238 0.00437597
R14178 VSS.n425 VSS.n424 0.00437597
R14179 VSS.n436 VSS.n435 0.00437597
R14180 VSS.n541 VSS.n540 0.00437597
R14181 VSS.n552 VSS.n544 0.00437597
R14182 VSS.n588 VSS.n587 0.00437597
R14183 VSS.n699 VSS.n698 0.00437597
R14184 VSS.n742 VSS.n741 0.00437597
R14185 VSS.n755 VSS.n745 0.00437597
R14186 VSS.n789 VSS.n788 0.00437597
R14187 VSS.n833 VSS.n832 0.00437597
R14188 VSS.n876 VSS.n875 0.00437597
R14189 VSS.n886 VSS.n879 0.00437597
R14190 VSS.n888 VSS.n691 0.0042037
R14191 VSS.n390 VSS.n389 0.00374675
R14192 VSS.n394 VSS.n393 0.00374675
R14193 VSS.n454 VSS.n453 0.00374675
R14194 VSS.n458 VSS.n457 0.00374675
R14195 VSS.n601 VSS.n600 0.00374675
R14196 VSS.n609 VSS.n608 0.00374675
R14197 VSS.n613 VSS.n612 0.00374675
R14198 VSS.n639 VSS.n638 0.00374675
R14199 VSS.n643 VSS.n642 0.00374675
R14200 VSS.n926 VSS.n925 0.00374675
R14201 VSS.n930 VSS.n929 0.00374675
R14202 VSS.n1080 VSS.n1079 0.00374675
R14203 VSS.n1084 VSS.n1083 0.00374675
R14204 VSS.n1256 VSS.n1255 0.00374675
R14205 VSS.n1260 VSS.n1259 0.00374675
R14206 VSS.n1404 VSS.n1403 0.00374675
R14207 VSS.n1408 VSS.n1407 0.00374675
R14208 VSS.n1548 VSS.n1547 0.00374675
R14209 VSS.n1552 VSS.n1551 0.00374675
R14210 VSS.n1697 VSS.n1693 0.00374675
R14211 VSS.n970 VSS.n961 0.00243798
R14212 VSS.n1147 VSS.n1140 0.00243798
R14213 VSS.n1300 VSS.n1290 0.00243798
R14214 VSS.n1450 VSS.n1443 0.00243798
R14215 VSS.n1599 VSS.n1582 0.00243798
R14216 VSS.n1667 VSS.n1666 0.00243798
R14217 VSS.n263 VSS.n262 0.00243798
R14218 VSS.n502 VSS.n495 0.00243798
R14219 VSS.n731 VSS.n721 0.00243798
R14220 VSS.n864 VSS.n855 0.00243798
R14221 VSS.n619 VSS.n618 0.00212338
R14222 VSS.n203 VSS.n202 0.00202439
R14223 VSS.n190 VSS.n189 0.00202439
R14224 VSS.n177 VSS.n176 0.00202439
R14225 VSS.n164 VSS.n163 0.00202439
R14226 VSS.n1025 VSS.n1024 0.00146899
R14227 VSS.n1180 VSS.n1179 0.00146899
R14228 VSS.n1333 VSS.n1332 0.00146899
R14229 VSS.n1495 VSS.n1494 0.00146899
R14230 VSS.n1636 VSS.n1635 0.00146899
R14231 VSS.n228 VSS.n209 0.00146899
R14232 VSS.n564 VSS.n563 0.00146899
R14233 VSS.n765 VSS.n764 0.00146899
R14234 VSS.n155 VSS.n154 0.000500344
R14235 pdrv2.n19 pdrv2.t177 92.4677
R14236 pdrv2.n19 pdrv2.t126 92.4677
R14237 pdrv2.n18 pdrv2.t81 92.4677
R14238 pdrv2.n18 pdrv2.t197 92.4677
R14239 pdrv2.n17 pdrv2.t146 92.4677
R14240 pdrv2.n17 pdrv2.t96 92.4677
R14241 pdrv2.n16 pdrv2.t55 92.4677
R14242 pdrv2.n16 pdrv2.t147 92.4677
R14243 pdrv2.n15 pdrv2.t50 92.4677
R14244 pdrv2.n15 pdrv2.t18 92.4677
R14245 pdrv2.n14 pdrv2.t165 92.4677
R14246 pdrv2.n14 pdrv2.t115 92.4677
R14247 pdrv2.n13 pdrv2.t70 92.4677
R14248 pdrv2.n13 pdrv2.t110 92.4677
R14249 pdrv2.n12 pdrv2.t64 92.4677
R14250 pdrv2.n12 pdrv2.t178 92.4677
R14251 pdrv2.n11 pdrv2.t187 92.4677
R14252 pdrv2.n11 pdrv2.t133 92.4677
R14253 pdrv2.n10 pdrv2.t44 92.4677
R14254 pdrv2.n10 pdrv2.t193 92.4677
R14255 pdrv2.n9 pdrv2.t86 92.4677
R14256 pdrv2.n9 pdrv2.t90 92.4677
R14257 pdrv2.n8 pdrv2.t13 92.4677
R14258 pdrv2.n8 pdrv2.t160 92.4677
R14259 pdrv2.n7 pdrv2.t112 92.4677
R14260 pdrv2.n7 pdrv2.t188 92.4677
R14261 pdrv2.n6 pdrv2.t42 92.4677
R14262 pdrv2.n6 pdrv2.t132 92.4677
R14263 pdrv2.n5 pdrv2.t186 92.4677
R14264 pdrv2.n5 pdrv2.t31 92.4677
R14265 pdrv2.n4 pdrv2.t116 92.4677
R14266 pdrv2.n4 pdrv2.t109 92.4677
R14267 pdrv2.n3 pdrv2.t10 92.4677
R14268 pdrv2.n3 pdrv2.t46 92.4677
R14269 pdrv2.n2 pdrv2.t139 92.4677
R14270 pdrv2.n2 pdrv2.t191 92.4677
R14271 pdrv2.n1 pdrv2.t184 92.4677
R14272 pdrv2.n1 pdrv2.t68 92.4677
R14273 pdrv2.n0 pdrv2.t190 92.4677
R14274 pdrv2.n0 pdrv2.t75 92.4677
R14275 pdrv2.n40 pdrv2.t102 92.465
R14276 pdrv2.n40 pdrv2.t21 92.465
R14277 pdrv2.n41 pdrv2.t91 92.465
R14278 pdrv2.n41 pdrv2.t11 92.465
R14279 pdrv2.n42 pdrv2.t22 92.465
R14280 pdrv2.n42 pdrv2.t168 92.465
R14281 pdrv2.n43 pdrv2.t66 92.465
R14282 pdrv2.n43 pdrv2.t32 92.465
R14283 pdrv2.n44 pdrv2.t136 92.465
R14284 pdrv2.n44 pdrv2.t145 92.465
R14285 pdrv2.n45 pdrv2.t49 92.465
R14286 pdrv2.n45 pdrv2.t16 92.465
R14287 pdrv2.n46 pdrv2.t162 92.465
R14288 pdrv2.n46 pdrv2.t62 92.465
R14289 pdrv2.n47 pdrv2.t20 92.465
R14290 pdrv2.n47 pdrv2.t138 92.465
R14291 pdrv2.n48 pdrv2.t189 92.465
R14292 pdrv2.n48 pdrv2.t33 92.465
R14293 pdrv2.n49 pdrv2.t118 92.465
R14294 pdrv2.n49 pdrv2.t113 92.465
R14295 pdrv2.n50 pdrv2.t23 92.465
R14296 pdrv2.n50 pdrv2.t63 92.465
R14297 pdrv2.n51 pdrv2.t163 92.465
R14298 pdrv2.n51 pdrv2.t17 92.465
R14299 pdrv2.n52 pdrv2.t9 92.465
R14300 pdrv2.n52 pdrv2.t89 92.465
R14301 pdrv2.n53 pdrv2.t137 92.465
R14302 pdrv2.n53 pdrv2.t95 92.465
R14303 pdrv2.n54 pdrv2.t144 92.465
R14304 pdrv2.n54 pdrv2.t195 92.465
R14305 pdrv2.n55 pdrv2.t37 92.465
R14306 pdrv2.n55 pdrv2.t73 92.465
R14307 pdrv2.n56 pdrv2.t175 92.465
R14308 pdrv2.n56 pdrv2.t80 92.465
R14309 pdrv2.n57 pdrv2.t124 92.465
R14310 pdrv2.n57 pdrv2.t174 92.465
R14311 pdrv2.n58 pdrv2.t27 92.465
R14312 pdrv2.n58 pdrv2.t107 92.465
R14313 pdrv2.n59 pdrv2.t158 92.465
R14314 pdrv2.n59 pdrv2.t5 92.465
R14315 pdrv2.n164 pdrv2.t12 92.4623
R14316 pdrv2.n165 pdrv2.t92 92.4623
R14317 pdrv2.n166 pdrv2.t141 92.4623
R14318 pdrv2.n167 pdrv2.t192 92.4623
R14319 pdrv2.n61 pdrv2.t65 92.4623
R14320 pdrv2.n61 pdrv2.t180 92.4623
R14321 pdrv2.n62 pdrv2.t57 92.4623
R14322 pdrv2.n62 pdrv2.t169 92.4623
R14323 pdrv2.n63 pdrv2.t181 92.4623
R14324 pdrv2.n63 pdrv2.t127 92.4623
R14325 pdrv2.n64 pdrv2.t38 92.4623
R14326 pdrv2.n64 pdrv2.t198 92.4623
R14327 pdrv2.n65 pdrv2.t97 92.4623
R14328 pdrv2.n65 pdrv2.t104 92.4623
R14329 pdrv2.n66 pdrv2.t24 92.4623
R14330 pdrv2.n66 pdrv2.t171 92.4623
R14331 pdrv2.n67 pdrv2.t119 92.4623
R14332 pdrv2.n67 pdrv2.t34 92.4623
R14333 pdrv2.n68 pdrv2.t179 92.4623
R14334 pdrv2.n68 pdrv2.t99 92.4623
R14335 pdrv2.n69 pdrv2.t149 92.4623
R14336 pdrv2.n69 pdrv2.t0 92.4623
R14337 pdrv2.n70 pdrv2.t83 92.4623
R14338 pdrv2.n70 pdrv2.t76 92.4623
R14339 pdrv2.n71 pdrv2.t182 92.4623
R14340 pdrv2.n71 pdrv2.t35 92.4623
R14341 pdrv2.n72 pdrv2.t122 92.4623
R14342 pdrv2.n72 pdrv2.t172 92.4623
R14343 pdrv2.n73 pdrv2.t166 92.4623
R14344 pdrv2.n73 pdrv2.t54 92.4623
R14345 pdrv2.n74 pdrv2.t98 92.4623
R14346 pdrv2.n74 pdrv2.t59 92.4623
R14347 pdrv2.n75 pdrv2.t103 92.4623
R14348 pdrv2.n75 pdrv2.t155 92.4623
R14349 pdrv2.n76 pdrv2.t3 92.4623
R14350 pdrv2.n76 pdrv2.t43 92.4623
R14351 pdrv2.n77 pdrv2.t131 92.4623
R14352 pdrv2.n77 pdrv2.t47 92.4623
R14353 pdrv2.n78 pdrv2.t85 92.4623
R14354 pdrv2.n78 pdrv2.t130 92.4623
R14355 pdrv2.n79 pdrv2.t185 92.4623
R14356 pdrv2.n79 pdrv2.t69 92.4623
R14357 pdrv2.n80 pdrv2.t114 92.4623
R14358 pdrv2.n80 pdrv2.t164 92.4623
R14359 pdrv2.n20 pdrv2.t45 92.4623
R14360 pdrv2.n20 pdrv2.t151 92.4623
R14361 pdrv2.n21 pdrv2.t39 92.4623
R14362 pdrv2.n21 pdrv2.t140 92.4623
R14363 pdrv2.n22 pdrv2.t150 92.4623
R14364 pdrv2.n22 pdrv2.t101 92.4623
R14365 pdrv2.n23 pdrv2.t19 92.4623
R14366 pdrv2.n23 pdrv2.t167 92.4623
R14367 pdrv2.n24 pdrv2.t71 92.4623
R14368 pdrv2.n24 pdrv2.t79 92.4623
R14369 pdrv2.n25 pdrv2.t196 92.4623
R14370 pdrv2.n25 pdrv2.t142 92.4623
R14371 pdrv2.n26 pdrv2.t93 92.4623
R14372 pdrv2.n26 pdrv2.t14 92.4623
R14373 pdrv2.n27 pdrv2.t148 92.4623
R14374 pdrv2.n27 pdrv2.t74 92.4623
R14375 pdrv2.n28 pdrv2.t117 92.4623
R14376 pdrv2.n28 pdrv2.t170 92.4623
R14377 pdrv2.n29 pdrv2.t58 92.4623
R14378 pdrv2.n29 pdrv2.t53 92.4623
R14379 pdrv2.n30 pdrv2.t154 92.4623
R14380 pdrv2.n30 pdrv2.t15 92.4623
R14381 pdrv2.n31 pdrv2.t94 92.4623
R14382 pdrv2.n31 pdrv2.t143 92.4623
R14383 pdrv2.n32 pdrv2.t135 92.4623
R14384 pdrv2.n32 pdrv2.t36 92.4623
R14385 pdrv2.n33 pdrv2.t72 92.4623
R14386 pdrv2.n33 pdrv2.t41 92.4623
R14387 pdrv2.n34 pdrv2.t78 92.4623
R14388 pdrv2.n34 pdrv2.t123 92.4623
R14389 pdrv2.n35 pdrv2.t173 92.4623
R14390 pdrv2.n35 pdrv2.t26 92.4623
R14391 pdrv2.n36 pdrv2.t106 92.4623
R14392 pdrv2.n36 pdrv2.t30 92.4623
R14393 pdrv2.n37 pdrv2.t61 92.4623
R14394 pdrv2.n37 pdrv2.t105 92.4623
R14395 pdrv2.n38 pdrv2.t157 92.4623
R14396 pdrv2.n38 pdrv2.t48 92.4623
R14397 pdrv2.n39 pdrv2.t88 92.4623
R14398 pdrv2.n39 pdrv2.t134 92.4623
R14399 pdrv2.n78 pdrv2.t159 92.4623
R14400 pdrv2.n78 pdrv2.t111 92.4623
R14401 pdrv2.n77 pdrv2.t67 92.4623
R14402 pdrv2.n77 pdrv2.t161 92.4623
R14403 pdrv2.n76 pdrv2.t60 92.4623
R14404 pdrv2.n76 pdrv2.t29 92.4623
R14405 pdrv2.n75 pdrv2.t183 92.4623
R14406 pdrv2.n75 pdrv2.t129 92.4623
R14407 pdrv2.n74 pdrv2.t84 92.4623
R14408 pdrv2.n74 pdrv2.t121 92.4623
R14409 pdrv2.n73 pdrv2.t77 92.4623
R14410 pdrv2.n73 pdrv2.t194 92.4623
R14411 pdrv2.n72 pdrv2.t2 92.4623
R14412 pdrv2.n72 pdrv2.t153 92.4623
R14413 pdrv2.n71 pdrv2.t52 92.4623
R14414 pdrv2.n71 pdrv2.t8 92.4623
R14415 pdrv2.n70 pdrv2.t100 92.4623
R14416 pdrv2.n70 pdrv2.t108 92.4623
R14417 pdrv2.n69 pdrv2.t28 92.4623
R14418 pdrv2.n69 pdrv2.t176 92.4623
R14419 pdrv2.n68 pdrv2.t125 92.4623
R14420 pdrv2.n68 pdrv2.t4 92.4623
R14421 pdrv2.n67 pdrv2.t51 92.4623
R14422 pdrv2.n67 pdrv2.t152 92.4623
R14423 pdrv2.n66 pdrv2.t1 92.4623
R14424 pdrv2.n66 pdrv2.t40 92.4623
R14425 pdrv2.n65 pdrv2.t128 92.4623
R14426 pdrv2.n65 pdrv2.t120 92.4623
R14427 pdrv2.n64 pdrv2.t25 92.4623
R14428 pdrv2.n64 pdrv2.t56 92.4623
R14429 pdrv2.n63 pdrv2.t156 92.4623
R14430 pdrv2.n63 pdrv2.t7 92.4623
R14431 pdrv2.n62 pdrv2.t199 92.4623
R14432 pdrv2.n62 pdrv2.t82 92.4623
R14433 pdrv2.n61 pdrv2.t6 92.4623
R14434 pdrv2.n61 pdrv2.t87 92.4623
R14435 pdrv2 pdrv2.n168 9.93689
R14436 pdrv2.n114 pdrv2.n113 1.02765
R14437 pdrv2.n124 pdrv2.n123 1.02179
R14438 pdrv2.n60 pdrv2.n132 0.989356
R14439 pdrv2.n126 pdrv2.n125 0.641125
R14440 pdrv2.n116 pdrv2.n115 0.641125
R14441 pdrv2.n133 pdrv2.n116 0.621594
R14442 pdrv2.n60 pdrv2.n126 0.621594
R14443 pdrv2.n115 pdrv2.n114 0.609875
R14444 pdrv2.n125 pdrv2.n124 0.609875
R14445 pdrv2.n168 pdrv2.n133 0.582531
R14446 pdrv2.n41 pdrv2.n40 0.515717
R14447 pdrv2.n21 pdrv2.n20 0.515717
R14448 pdrv2.n1 pdrv2.n0 0.515717
R14449 pdrv2.n168 pdrv2.n167 0.398889
R14450 pdrv2.n61 pdrv2.n60 0.396152
R14451 pdrv2.n80 pdrv2.n79 0.343978
R14452 pdrv2.n79 pdrv2.n78 0.343978
R14453 pdrv2.n78 pdrv2.n77 0.343978
R14454 pdrv2.n77 pdrv2.n76 0.343978
R14455 pdrv2.n76 pdrv2.n75 0.343978
R14456 pdrv2.n75 pdrv2.n74 0.343978
R14457 pdrv2.n74 pdrv2.n73 0.343978
R14458 pdrv2.n73 pdrv2.n72 0.343978
R14459 pdrv2.n72 pdrv2.n71 0.343978
R14460 pdrv2.n71 pdrv2.n70 0.343978
R14461 pdrv2.n70 pdrv2.n69 0.343978
R14462 pdrv2.n69 pdrv2.n68 0.343978
R14463 pdrv2.n68 pdrv2.n67 0.343978
R14464 pdrv2.n67 pdrv2.n66 0.343978
R14465 pdrv2.n66 pdrv2.n65 0.343978
R14466 pdrv2.n65 pdrv2.n64 0.343978
R14467 pdrv2.n64 pdrv2.n63 0.343978
R14468 pdrv2.n63 pdrv2.n62 0.343978
R14469 pdrv2.n62 pdrv2.n61 0.343978
R14470 pdrv2.n59 pdrv2.n58 0.343978
R14471 pdrv2.n58 pdrv2.n57 0.343978
R14472 pdrv2.n57 pdrv2.n56 0.343978
R14473 pdrv2.n56 pdrv2.n55 0.343978
R14474 pdrv2.n55 pdrv2.n54 0.343978
R14475 pdrv2.n54 pdrv2.n53 0.343978
R14476 pdrv2.n53 pdrv2.n52 0.343978
R14477 pdrv2.n52 pdrv2.n51 0.343978
R14478 pdrv2.n51 pdrv2.n50 0.343978
R14479 pdrv2.n50 pdrv2.n49 0.343978
R14480 pdrv2.n49 pdrv2.n48 0.343978
R14481 pdrv2.n48 pdrv2.n47 0.343978
R14482 pdrv2.n47 pdrv2.n46 0.343978
R14483 pdrv2.n46 pdrv2.n45 0.343978
R14484 pdrv2.n45 pdrv2.n44 0.343978
R14485 pdrv2.n44 pdrv2.n43 0.343978
R14486 pdrv2.n43 pdrv2.n42 0.343978
R14487 pdrv2.n42 pdrv2.n41 0.343978
R14488 pdrv2.n39 pdrv2.n38 0.343978
R14489 pdrv2.n38 pdrv2.n37 0.343978
R14490 pdrv2.n37 pdrv2.n36 0.343978
R14491 pdrv2.n36 pdrv2.n35 0.343978
R14492 pdrv2.n35 pdrv2.n34 0.343978
R14493 pdrv2.n34 pdrv2.n33 0.343978
R14494 pdrv2.n33 pdrv2.n32 0.343978
R14495 pdrv2.n32 pdrv2.n31 0.343978
R14496 pdrv2.n31 pdrv2.n30 0.343978
R14497 pdrv2.n30 pdrv2.n29 0.343978
R14498 pdrv2.n29 pdrv2.n28 0.343978
R14499 pdrv2.n28 pdrv2.n27 0.343978
R14500 pdrv2.n27 pdrv2.n26 0.343978
R14501 pdrv2.n26 pdrv2.n25 0.343978
R14502 pdrv2.n25 pdrv2.n24 0.343978
R14503 pdrv2.n24 pdrv2.n23 0.343978
R14504 pdrv2.n23 pdrv2.n22 0.343978
R14505 pdrv2.n22 pdrv2.n21 0.343978
R14506 pdrv2.n19 pdrv2.n18 0.343978
R14507 pdrv2.n18 pdrv2.n17 0.343978
R14508 pdrv2.n17 pdrv2.n16 0.343978
R14509 pdrv2.n16 pdrv2.n15 0.343978
R14510 pdrv2.n15 pdrv2.n14 0.343978
R14511 pdrv2.n14 pdrv2.n13 0.343978
R14512 pdrv2.n13 pdrv2.n12 0.343978
R14513 pdrv2.n12 pdrv2.n11 0.343978
R14514 pdrv2.n11 pdrv2.n10 0.343978
R14515 pdrv2.n10 pdrv2.n9 0.343978
R14516 pdrv2.n9 pdrv2.n8 0.343978
R14517 pdrv2.n8 pdrv2.n7 0.343978
R14518 pdrv2.n7 pdrv2.n6 0.343978
R14519 pdrv2.n6 pdrv2.n5 0.343978
R14520 pdrv2.n5 pdrv2.n4 0.343978
R14521 pdrv2.n4 pdrv2.n3 0.343978
R14522 pdrv2.n3 pdrv2.n2 0.343978
R14523 pdrv2.n2 pdrv2.n1 0.343978
R14524 pdrv2.n167 pdrv2.n166 0.298524
R14525 pdrv2.n166 pdrv2.n165 0.298524
R14526 pdrv2.n165 pdrv2.n164 0.298524
R14527 pdrv2.n164 pdrv2.n163 0.298524
R14528 pdrv2.n163 pdrv2.n162 0.298524
R14529 pdrv2.n162 pdrv2.n161 0.298524
R14530 pdrv2.n161 pdrv2.n160 0.298524
R14531 pdrv2.n160 pdrv2.n159 0.298524
R14532 pdrv2.n159 pdrv2.n158 0.298524
R14533 pdrv2.n158 pdrv2.n157 0.298524
R14534 pdrv2.n157 pdrv2.n156 0.298524
R14535 pdrv2.n156 pdrv2.n155 0.298524
R14536 pdrv2.n155 pdrv2.n154 0.298524
R14537 pdrv2.n154 pdrv2.n153 0.298524
R14538 pdrv2.n153 pdrv2.n152 0.298524
R14539 pdrv2.n152 pdrv2.n151 0.298524
R14540 pdrv2.n151 pdrv2.n150 0.298524
R14541 pdrv2.n150 pdrv2.n149 0.298524
R14542 pdrv2.n149 pdrv2.n148 0.298524
R14543 pdrv2.n148 pdrv2.n147 0.298524
R14544 pdrv2.n147 pdrv2.n146 0.298524
R14545 pdrv2.n146 pdrv2.n145 0.298524
R14546 pdrv2.n145 pdrv2.n144 0.298524
R14547 pdrv2.n144 pdrv2.n143 0.298524
R14548 pdrv2.n143 pdrv2.n142 0.298524
R14549 pdrv2.n142 pdrv2.n141 0.298524
R14550 pdrv2.n141 pdrv2.n140 0.298524
R14551 pdrv2.n140 pdrv2.n139 0.298524
R14552 pdrv2.n139 pdrv2.n138 0.298524
R14553 pdrv2.n138 pdrv2.n137 0.298524
R14554 pdrv2.n137 pdrv2.n136 0.298524
R14555 pdrv2.n136 pdrv2.n135 0.298524
R14556 pdrv2.n135 pdrv2.n134 0.298524
R14557 pdrv2.n128 pdrv2.n127 0.298524
R14558 pdrv2.n129 pdrv2.n128 0.298524
R14559 pdrv2.n130 pdrv2.n129 0.298524
R14560 pdrv2.n131 pdrv2.n130 0.298524
R14561 pdrv2.n132 pdrv2.n131 0.298524
R14562 pdrv2.n123 pdrv2.n122 0.26965
R14563 pdrv2.n122 pdrv2.n121 0.26965
R14564 pdrv2.n121 pdrv2.n120 0.26965
R14565 pdrv2.n120 pdrv2.n119 0.26965
R14566 pdrv2.n119 pdrv2.n118 0.26965
R14567 pdrv2.n118 pdrv2.n117 0.26965
R14568 pdrv2.n82 pdrv2.n81 0.26965
R14569 pdrv2.n83 pdrv2.n82 0.26965
R14570 pdrv2.n84 pdrv2.n83 0.26965
R14571 pdrv2.n85 pdrv2.n84 0.26965
R14572 pdrv2.n86 pdrv2.n85 0.26965
R14573 pdrv2.n87 pdrv2.n86 0.26965
R14574 pdrv2.n88 pdrv2.n87 0.26965
R14575 pdrv2.n89 pdrv2.n88 0.26965
R14576 pdrv2.n90 pdrv2.n89 0.26965
R14577 pdrv2.n91 pdrv2.n90 0.26965
R14578 pdrv2.n92 pdrv2.n91 0.26965
R14579 pdrv2.n93 pdrv2.n92 0.26965
R14580 pdrv2.n94 pdrv2.n93 0.26965
R14581 pdrv2.n95 pdrv2.n94 0.26965
R14582 pdrv2.n96 pdrv2.n95 0.26965
R14583 pdrv2.n97 pdrv2.n96 0.26965
R14584 pdrv2.n98 pdrv2.n97 0.26965
R14585 pdrv2.n99 pdrv2.n98 0.26965
R14586 pdrv2.n100 pdrv2.n99 0.26965
R14587 pdrv2.n101 pdrv2.n100 0.26965
R14588 pdrv2.n102 pdrv2.n101 0.26965
R14589 pdrv2.n103 pdrv2.n102 0.26965
R14590 pdrv2.n104 pdrv2.n103 0.26965
R14591 pdrv2.n105 pdrv2.n104 0.26965
R14592 pdrv2.n106 pdrv2.n105 0.26965
R14593 pdrv2.n107 pdrv2.n106 0.26965
R14594 pdrv2.n108 pdrv2.n107 0.26965
R14595 pdrv2.n109 pdrv2.n108 0.26965
R14596 pdrv2.n110 pdrv2.n109 0.26965
R14597 pdrv2.n111 pdrv2.n110 0.26965
R14598 pdrv2.n112 pdrv2.n111 0.26965
R14599 pdrv2.n113 pdrv2.n112 0.26965
R14600 pdrv2.n114 pdrv2.n19 0.227674
R14601 pdrv2.n115 pdrv2.n39 0.227674
R14602 pdrv2.n116 pdrv2.n59 0.227674
R14603 pdrv2.n133 pdrv2.n80 0.227674
R14604 nbias.n7 nbias.t4 88.61
R14605 nbias.n2 nbias.t10 88.1243
R14606 nbias.n7 nbias.t0 88.1243
R14607 nbias.n8 nbias.t6 88.1243
R14608 nbias.n9 nbias.t2 88.1243
R14609 nbias.n15 nbias.t9 50.3368
R14610 nbias.n15 nbias.t11 46.6005
R14611 nbias.n3 nbias.t8 23.2945
R14612 nbias.n16 nbias.t1 16.5305
R14613 nbias.n16 nbias.t5 16.5305
R14614 nbias.n23 nbias.t3 16.5305
R14615 nbias.n23 nbias.t7 16.5305
R14616 nbias.n0 nbias.n18 9.32489
R14617 nbias.n1 nbias.n25 9.32489
R14618 nbias.n17 nbias.n16 8.35
R14619 nbias.n24 nbias.n23 8.34928
R14620 nbias.n0 nbias.n20 4.5005
R14621 nbias.n1 nbias.n27 4.5005
R14622 nbias.n22 nbias.n15 3.93502
R14623 nbias.n0 nbias.n17 2.34459
R14624 nbias.n1 nbias.n24 2.34448
R14625 nbias.n30 nbias.n14 1.39011
R14626 nbias.n28 nbias.n1 0.88838
R14627 nbias.n21 nbias.n0 0.888379
R14628 nbias.n4 nbias.n3 0.87589
R14629 nbias.n14 nbias.n9 0.871132
R14630 nbias.n3 nbias.n2 0.863003
R14631 nbias nbias.n30 0.771333
R14632 nbias.n13 nbias.n12 0.717167
R14633 nbias.n29 nbias.n22 0.690976
R14634 nbias.n30 nbias.n29 0.664191
R14635 nbias.n12 nbias.n11 0.5255
R14636 nbias.n11 nbias.n10 0.5255
R14637 nbias.n8 nbias.n7 0.486214
R14638 nbias.n9 nbias.n8 0.486214
R14639 nbias.n20 nbias.n19 0.376971
R14640 nbias.n27 nbias.n26 0.376971
R14641 nbias nbias.n6 0.278669
R14642 nbias.n22 nbias.n21 0.243398
R14643 nbias.n29 nbias.n28 0.243398
R14644 nbias.n14 nbias.n13 0.219013
R14645 nbias.n6 nbias.n5 0.113176
R14646 nbias.n5 nbias.n4 0.113176
R14647 VIN.n0 VIN.t2 93.5207
R14648 VIN.n0 VIN.t3 93.5037
R14649 VIN.n2 VIN.t0 46.1462
R14650 VIN.n1 VIN.t1 46.105
R14651 VIN.n1 VIN.n0 5.25741
R14652 VIN.n2 VIN.n1 3.166
R14653 VIN VIN.n2 0.59831
R14654 EN.n0 EN.t1 63.176
R14655 EN.n0 EN.t0 5.00531
R14656 EN EN.n0 0.717948
R14657 VIP.n0 VIP.t3 93.2353
R14658 VIP.n0 VIP.t0 93.2134
R14659 VIP.n1 VIP.t2 46.4551
R14660 VIP.n2 VIP.t1 46.4185
R14661 VIP VIP.n2 3.37627
R14662 VIP.n2 VIP.n1 3.23285
R14663 VIP.n1 VIP.n0 2.72991
C0 pbias VOUT 0.00123f
C1 nbias VDD 0.0967f
C2 vcomn2 VSS 0.674f
C3 vcomp a_n551_n345# 0.51f
C4 VOUT VIN 0.00329f
C5 VSS EN 1.77f
C6 a_n1922_640# EN 0.0495f
C7 a_n3090_640# VDD 2f
C8 pdrv2 VOUT 32.6f
C9 pdrv1 VSS 0.879f
C10 pdrv1 a_n1922_640# 0.506f
C11 a_1610_n2436# a_1610_n3072# 0.141f
C12 nbias VSS 5.38f
C13 vcomn1 VDD 0.0047f
C14 ndrv VDD 0.923f
C15 a_n1922_640# nbias 0.0546f
C16 VOUT EN 0.00603f
C17 VIP VIN 1.54f
C18 a_n3822_n2754# a_n3822_n3390# 0.14f
C19 pdrv1 VOUT 31.9f
C20 pdrv2 VIP 1.24f
C21 a_n3090_640# VSS 0.358f
C22 a_n3090_640# a_n1922_640# 0.00662f
C23 vcomn1 VSS 0.593f
C24 a_1610_n2436# VDD 1.77f
C25 vcomn2 VIP 0.233f
C26 pbias VIN 0.0456f
C27 nbias VOUT 0.0229f
C28 vcomp VDD 1.35f
C29 ndrv VSS 45.8f
C30 a_n1922_640# vcomn1 0.214f
C31 VIP EN 0.31f
C32 a_n1922_640# ndrv 0.0061f
C33 a_n3090_640# VOUT 2.79e-19
C34 pdrv2 VIN 0.0733f
C35 pdrv1 VIP 0.858f
C36 vcomn2 VIN 0.231f
C37 pbias EN 0.0456f
C38 nbias VIP 0.0624f
C39 a_1610_n2436# VSS 1.61f
C40 vcomp VSS 0.00513f
C41 a_n551_n345# VDD 0.423f
C42 ndrv VOUT 19.1f
C43 VIN EN 2.17f
C44 a_n1922_640# vcomp 0.00829f
C45 pdrv1 pbias 0.139f
C46 pdrv2 vcomn2 0.181f
C47 a_n3090_640# VIP 0.203f
C48 pdrv1 VIN 0.546f
C49 pdrv2 EN 0.0663f
C50 pdrv2 pdrv1 1.46f
C51 a_1610_n3072# VDD 0.194f
C52 pbias nbias 0.344f
C53 ndrv a_n3822_n2754# 0.00331f
C54 nbias VIN 0.0903f
C55 a_1610_n2436# VOUT 0.651f
C56 vcomn1 VIP 0.228f
C57 vcomn2 EN 0.187f
C58 ndrv VIP 0.396f
C59 a_n551_n345# VSS 1.73f
C60 pdrv2 nbias 0.0365f
C61 pdrv1 EN 0.144f
C62 a_n3090_640# VIN 0.336f
C63 pdrv2 a_n3090_640# 0.714f
C64 a_1610_n3072# VSS 0.316f
C65 vcomn2 nbias 0.284f
C66 ndrv pbias 0.00129f
C67 vcomn1 VIN 0.233f
C68 nbias EN 1.81f
C69 ndrv VIN 0.125f
C70 a_n551_n345# VOUT 4.88e-19
C71 vcomp VIP 0.145f
C72 a_n3090_640# vcomn2 0.226f
C73 pdrv1 nbias 0.0901f
C74 pdrv2 ndrv 0.00332f
C75 a_n3090_640# EN 0.0688f
C76 ndrv a_n3822_n3390# 7.3e-19
C77 pdrv1 a_n3090_640# 0.0067f
C78 vcomn2 vcomn1 0.0723f
C79 ndrv vcomn2 0.266f
C80 vcomp pbias 0.162f
C81 vcomn1 EN 0.00189f
C82 VDD VSS 0.109p
C83 a_n551_n345# VIP 0.00414f
C84 ndrv EN 0.206f
C85 vcomp VIN 0.144f
C86 a_n1922_640# VDD 1.94f
C87 pdrv1 vcomn1 0.17f
C88 a_n3090_640# nbias 0.00341f
C89 pdrv1 ndrv 0.209f
C90 pdrv2 vcomp 1.65e-19
C91 nbias vcomn1 0.601f
C92 a_n551_n345# pbias 0.0349f
C93 ndrv nbias 0.296f
C94 a_1610_n2436# EN 0.151f
C95 VDD VOUT 0.12p
C96 a_n551_n345# VIN 0.506f
C97 vcomp EN 1.78e-19
C98 a_n1922_640# VSS 0.341f
C99 pdrv1 a_1610_n2436# 0.0145f
C100 pdrv1 vcomp 0.398f
C101 a_n3090_640# ndrv 0.0064f
C102 nbias a_1610_n2436# 0.0399f
C103 ndrv vcomn1 0.324f
C104 vcomp nbias 0.00684f
C105 VDD VIP 1.27f
C106 VSS VOUT 34.6f
C107 a_n551_n345# EN 0.154f
C108 a_n1922_640# VOUT 4.05e-19
C109 pdrv1 a_n551_n345# 0.0987f
C110 a_n3090_640# vcomp 4.79e-19
C111 a_n3822_n2754# VSS 0.58f
C112 pbias VDD 1.29f
C113 ndrv a_1610_n2436# 0.635f
C114 a_n551_n345# nbias 0.311f
C115 ndrv vcomp 0.427f
C116 VDD VIN 0.609f
C117 VSS VIP 1.45f
C118 a_n1922_640# VIP 0.224f
C119 pdrv2 VDD 71.2f
C120 pbias VSS 0.4f
C121 vcomn2 VDD 5.13e-19
C122 a_n551_n345# vcomn1 0.00534f
C123 ndrv a_n551_n345# 0.465f
C124 VSS VIN 1.17f
C125 VOUT VIP 3.71e-19
C126 VDD EN 0.311f
C127 a_n1922_640# VIN 0.36f
C128 pdrv2 VSS 0.699f
C129 pdrv1 VDD 67.9f
C130 pdrv2 a_n1922_640# 0.0981f
C131 a_n3822_n3390# VSS 0.563f
C132 ndrv a_1610_n3072# 0.0012f
C133 EN VSUBS 0.448f
C134 VIN VSUBS 0.357f
C135 VIP VSUBS 0.407f
C136 VOUT VSUBS 7.09f
C137 VSS VSUBS 0.739f
C138 VDD VSUBS 0.239p
C139 a_n3822_n3390# VSUBS 0.393f
C140 a_1610_n3072# VSUBS 0.413f
C141 a_n3822_n2754# VSUBS 0.379f
C142 a_1610_n2436# VSUBS 0.213f
C143 vcomn1 VSUBS 0.0488f
C144 nbias VSUBS 0.535f
C145 vcomn2 VSUBS 0.0488f
C146 pbias VSUBS 0.212f
C147 a_n551_n345# VSUBS 0.177f
C148 vcomp VSUBS 0.0721f
C149 ndrv VSUBS 11.2f
C150 a_n1922_640# VSUBS 0.287f
C151 a_n3090_640# VSUBS 0.288f
C152 pdrv1 VSUBS 13.8f
C153 pdrv2 VSUBS 16.2f
C154 EN.t0 VSUBS 0.136f
C155 EN.t1 VSUBS 0.339f
C156 EN.n0 VSUBS 1.43f
C157 VIN.t2 VSUBS 0.1f
C158 VIN.t3 VSUBS 0.1f
C159 VIN.n0 VSUBS 0.364f
C160 VIN.t1 VSUBS 0.123f
C161 VIN.n1 VSUBS 0.776f
C162 VIN.t0 VSUBS 0.123f
C163 VIN.n2 VSUBS 0.559f
C164 nbias.n0 VSUBS 0.102f
C165 nbias.n1 VSUBS 0.102f
C166 nbias.t10 VSUBS 0.121f
C167 nbias.n2 VSUBS 0.132f
C168 nbias.t8 VSUBS 0.0407f
C169 nbias.n3 VSUBS 0.501f
C170 nbias.n4 VSUBS 0.103f
C171 nbias.n5 VSUBS 0.0284f
C172 nbias.n6 VSUBS 0.0431f
C173 nbias.t2 VSUBS 0.12f
C174 nbias.t6 VSUBS 0.12f
C175 nbias.t0 VSUBS 0.12f
C176 nbias.t4 VSUBS 0.121f
C177 nbias.n7 VSUBS 0.231f
C178 nbias.n8 VSUBS 0.12f
C179 nbias.n9 VSUBS 0.144f
C180 nbias.n10 VSUBS 0.228f
C181 nbias.n11 VSUBS 0.118f
C182 nbias.n12 VSUBS 0.121f
C183 nbias.n13 VSUBS 0.0823f
C184 nbias.n14 VSUBS 0.168f
C185 nbias.t11 VSUBS 0.137f
C186 nbias.t9 VSUBS 0.174f
C187 nbias.n15 VSUBS 1.11f
C188 nbias.t1 VSUBS 0.0181f
C189 nbias.t5 VSUBS 0.0181f
C190 nbias.n16 VSUBS 0.0399f
C191 nbias.n17 VSUBS 0.0111f
C192 nbias.n18 VSUBS 0.0122f
C193 nbias.n19 VSUBS 0.00753f
C194 nbias.n20 VSUBS 0.00181f
C195 nbias.n21 VSUBS 0.109f
C196 nbias.n22 VSUBS 0.263f
C197 nbias.t3 VSUBS 0.0181f
C198 nbias.t7 VSUBS 0.0181f
C199 nbias.n23 VSUBS 0.0399f
C200 nbias.n24 VSUBS 0.0111f
C201 nbias.n25 VSUBS 0.0122f
C202 nbias.n26 VSUBS 0.00753f
C203 nbias.n27 VSUBS 0.00181f
C204 nbias.n28 VSUBS 0.109f
C205 nbias.n29 VSUBS 0.118f
C206 nbias.n30 VSUBS 0.248f
C207 pdrv2.n0 VSUBS 0.707f
C208 pdrv2.n1 VSUBS 0.686f
C209 pdrv2.n2 VSUBS 0.686f
C210 pdrv2.n3 VSUBS 0.686f
C211 pdrv2.n4 VSUBS 0.686f
C212 pdrv2.n5 VSUBS 0.686f
C213 pdrv2.n6 VSUBS 0.686f
C214 pdrv2.n7 VSUBS 0.686f
C215 pdrv2.n8 VSUBS 0.686f
C216 pdrv2.n9 VSUBS 0.686f
C217 pdrv2.n10 VSUBS 0.686f
C218 pdrv2.n11 VSUBS 0.686f
C219 pdrv2.n12 VSUBS 0.686f
C220 pdrv2.n13 VSUBS 0.686f
C221 pdrv2.n14 VSUBS 0.686f
C222 pdrv2.n15 VSUBS 0.686f
C223 pdrv2.n16 VSUBS 0.686f
C224 pdrv2.n17 VSUBS 0.686f
C225 pdrv2.n18 VSUBS 0.686f
C226 pdrv2.n19 VSUBS 0.708f
C227 pdrv2.n20 VSUBS 0.633f
C228 pdrv2.n21 VSUBS 0.612f
C229 pdrv2.n22 VSUBS 0.612f
C230 pdrv2.n23 VSUBS 0.612f
C231 pdrv2.n24 VSUBS 0.612f
C232 pdrv2.n25 VSUBS 0.612f
C233 pdrv2.n26 VSUBS 0.612f
C234 pdrv2.n27 VSUBS 0.612f
C235 pdrv2.n28 VSUBS 0.612f
C236 pdrv2.n29 VSUBS 0.612f
C237 pdrv2.n30 VSUBS 0.612f
C238 pdrv2.n31 VSUBS 0.612f
C239 pdrv2.n32 VSUBS 0.612f
C240 pdrv2.n33 VSUBS 0.612f
C241 pdrv2.n34 VSUBS 0.612f
C242 pdrv2.n35 VSUBS 0.612f
C243 pdrv2.n36 VSUBS 0.612f
C244 pdrv2.n37 VSUBS 0.612f
C245 pdrv2.n38 VSUBS 0.612f
C246 pdrv2.n39 VSUBS 0.634f
C247 pdrv2.n40 VSUBS 0.702f
C248 pdrv2.n41 VSUBS 0.681f
C249 pdrv2.n42 VSUBS 0.681f
C250 pdrv2.n43 VSUBS 0.681f
C251 pdrv2.n44 VSUBS 0.681f
C252 pdrv2.n45 VSUBS 0.681f
C253 pdrv2.n46 VSUBS 0.681f
C254 pdrv2.n47 VSUBS 0.681f
C255 pdrv2.n48 VSUBS 0.681f
C256 pdrv2.n49 VSUBS 0.681f
C257 pdrv2.n50 VSUBS 0.681f
C258 pdrv2.n51 VSUBS 0.681f
C259 pdrv2.n52 VSUBS 0.681f
C260 pdrv2.n53 VSUBS 0.681f
C261 pdrv2.n54 VSUBS 0.681f
C262 pdrv2.n55 VSUBS 0.681f
C263 pdrv2.n56 VSUBS 0.681f
C264 pdrv2.n57 VSUBS 0.681f
C265 pdrv2.n58 VSUBS 0.681f
C266 pdrv2.n59 VSUBS 0.703f
C267 pdrv2.n60 VSUBS 0.321f
C268 pdrv2.n61 VSUBS 0.633f
C269 pdrv2.n62 VSUBS 0.612f
C270 pdrv2.n63 VSUBS 0.612f
C271 pdrv2.n64 VSUBS 0.612f
C272 pdrv2.n65 VSUBS 0.612f
C273 pdrv2.n66 VSUBS 0.612f
C274 pdrv2.n67 VSUBS 0.612f
C275 pdrv2.n68 VSUBS 0.612f
C276 pdrv2.n69 VSUBS 0.612f
C277 pdrv2.n70 VSUBS 0.612f
C278 pdrv2.n71 VSUBS 0.612f
C279 pdrv2.n72 VSUBS 0.612f
C280 pdrv2.n73 VSUBS 0.612f
C281 pdrv2.n74 VSUBS 0.612f
C282 pdrv2.n75 VSUBS 0.612f
C283 pdrv2.n76 VSUBS 0.612f
C284 pdrv2.n77 VSUBS 0.612f
C285 pdrv2.n78 VSUBS 0.612f
C286 pdrv2.n79 VSUBS 0.612f
C287 pdrv2.n80 VSUBS 0.634f
C288 pdrv2.n81 VSUBS 0.187f
C289 pdrv2.n82 VSUBS 0.187f
C290 pdrv2.n83 VSUBS 0.187f
C291 pdrv2.n84 VSUBS 0.187f
C292 pdrv2.n85 VSUBS 0.187f
C293 pdrv2.n86 VSUBS 0.187f
C294 pdrv2.n87 VSUBS 0.187f
C295 pdrv2.n88 VSUBS 0.187f
C296 pdrv2.n89 VSUBS 0.187f
C297 pdrv2.n90 VSUBS 0.187f
C298 pdrv2.n91 VSUBS 0.187f
C299 pdrv2.n92 VSUBS 0.187f
C300 pdrv2.n93 VSUBS 0.187f
C301 pdrv2.n94 VSUBS 0.187f
C302 pdrv2.n95 VSUBS 0.187f
C303 pdrv2.n96 VSUBS 0.187f
C304 pdrv2.n97 VSUBS 0.187f
C305 pdrv2.n98 VSUBS 0.187f
C306 pdrv2.n99 VSUBS 0.187f
C307 pdrv2.n100 VSUBS 0.187f
C308 pdrv2.n101 VSUBS 0.187f
C309 pdrv2.n102 VSUBS 0.187f
C310 pdrv2.n103 VSUBS 0.187f
C311 pdrv2.n104 VSUBS 0.187f
C312 pdrv2.n105 VSUBS 0.187f
C313 pdrv2.n106 VSUBS 0.187f
C314 pdrv2.n107 VSUBS 0.187f
C315 pdrv2.n108 VSUBS 0.187f
C316 pdrv2.n109 VSUBS 0.187f
C317 pdrv2.n110 VSUBS 0.187f
C318 pdrv2.n111 VSUBS 0.187f
C319 pdrv2.n112 VSUBS 0.187f
C320 pdrv2.n113 VSUBS 0.289f
C321 pdrv2.t177 VSUBS 0.151f
C322 pdrv2.t126 VSUBS 0.151f
C323 pdrv2.t81 VSUBS 0.151f
C324 pdrv2.t197 VSUBS 0.151f
C325 pdrv2.t146 VSUBS 0.151f
C326 pdrv2.t96 VSUBS 0.151f
C327 pdrv2.t55 VSUBS 0.151f
C328 pdrv2.t147 VSUBS 0.151f
C329 pdrv2.t50 VSUBS 0.151f
C330 pdrv2.t18 VSUBS 0.151f
C331 pdrv2.t165 VSUBS 0.151f
C332 pdrv2.t115 VSUBS 0.151f
C333 pdrv2.t70 VSUBS 0.151f
C334 pdrv2.t110 VSUBS 0.151f
C335 pdrv2.t64 VSUBS 0.151f
C336 pdrv2.t178 VSUBS 0.151f
C337 pdrv2.t187 VSUBS 0.151f
C338 pdrv2.t133 VSUBS 0.151f
C339 pdrv2.t44 VSUBS 0.151f
C340 pdrv2.t193 VSUBS 0.151f
C341 pdrv2.t86 VSUBS 0.151f
C342 pdrv2.t90 VSUBS 0.151f
C343 pdrv2.t13 VSUBS 0.151f
C344 pdrv2.t160 VSUBS 0.151f
C345 pdrv2.t112 VSUBS 0.151f
C346 pdrv2.t188 VSUBS 0.151f
C347 pdrv2.t42 VSUBS 0.151f
C348 pdrv2.t132 VSUBS 0.151f
C349 pdrv2.t186 VSUBS 0.151f
C350 pdrv2.t31 VSUBS 0.151f
C351 pdrv2.t116 VSUBS 0.151f
C352 pdrv2.t109 VSUBS 0.151f
C353 pdrv2.t10 VSUBS 0.151f
C354 pdrv2.t46 VSUBS 0.151f
C355 pdrv2.t139 VSUBS 0.151f
C356 pdrv2.t191 VSUBS 0.151f
C357 pdrv2.t184 VSUBS 0.151f
C358 pdrv2.t68 VSUBS 0.151f
C359 pdrv2.t190 VSUBS 0.151f
C360 pdrv2.t75 VSUBS 0.151f
C361 pdrv2.n114 VSUBS 0.326f
C362 pdrv2.t45 VSUBS 0.151f
C363 pdrv2.t151 VSUBS 0.151f
C364 pdrv2.t39 VSUBS 0.151f
C365 pdrv2.t140 VSUBS 0.151f
C366 pdrv2.t150 VSUBS 0.151f
C367 pdrv2.t101 VSUBS 0.151f
C368 pdrv2.t19 VSUBS 0.151f
C369 pdrv2.t167 VSUBS 0.151f
C370 pdrv2.t71 VSUBS 0.151f
C371 pdrv2.t79 VSUBS 0.151f
C372 pdrv2.t196 VSUBS 0.151f
C373 pdrv2.t142 VSUBS 0.151f
C374 pdrv2.t93 VSUBS 0.151f
C375 pdrv2.t14 VSUBS 0.151f
C376 pdrv2.t148 VSUBS 0.151f
C377 pdrv2.t74 VSUBS 0.151f
C378 pdrv2.t117 VSUBS 0.151f
C379 pdrv2.t170 VSUBS 0.151f
C380 pdrv2.t58 VSUBS 0.151f
C381 pdrv2.t53 VSUBS 0.151f
C382 pdrv2.t154 VSUBS 0.151f
C383 pdrv2.t15 VSUBS 0.151f
C384 pdrv2.t94 VSUBS 0.151f
C385 pdrv2.t143 VSUBS 0.151f
C386 pdrv2.t135 VSUBS 0.151f
C387 pdrv2.t36 VSUBS 0.151f
C388 pdrv2.t72 VSUBS 0.151f
C389 pdrv2.t41 VSUBS 0.151f
C390 pdrv2.t78 VSUBS 0.151f
C391 pdrv2.t123 VSUBS 0.151f
C392 pdrv2.t173 VSUBS 0.151f
C393 pdrv2.t26 VSUBS 0.151f
C394 pdrv2.t106 VSUBS 0.151f
C395 pdrv2.t30 VSUBS 0.151f
C396 pdrv2.t61 VSUBS 0.151f
C397 pdrv2.t105 VSUBS 0.151f
C398 pdrv2.t157 VSUBS 0.151f
C399 pdrv2.t48 VSUBS 0.151f
C400 pdrv2.t88 VSUBS 0.151f
C401 pdrv2.t134 VSUBS 0.151f
C402 pdrv2.n115 VSUBS 0.272f
C403 pdrv2.t5 VSUBS 0.151f
C404 pdrv2.t158 VSUBS 0.151f
C405 pdrv2.t107 VSUBS 0.151f
C406 pdrv2.t27 VSUBS 0.151f
C407 pdrv2.t174 VSUBS 0.151f
C408 pdrv2.t124 VSUBS 0.151f
C409 pdrv2.t80 VSUBS 0.151f
C410 pdrv2.t175 VSUBS 0.151f
C411 pdrv2.t73 VSUBS 0.151f
C412 pdrv2.t37 VSUBS 0.151f
C413 pdrv2.t195 VSUBS 0.151f
C414 pdrv2.t144 VSUBS 0.151f
C415 pdrv2.t95 VSUBS 0.151f
C416 pdrv2.t137 VSUBS 0.151f
C417 pdrv2.t89 VSUBS 0.151f
C418 pdrv2.t9 VSUBS 0.151f
C419 pdrv2.t17 VSUBS 0.151f
C420 pdrv2.t163 VSUBS 0.151f
C421 pdrv2.t63 VSUBS 0.151f
C422 pdrv2.t23 VSUBS 0.151f
C423 pdrv2.t113 VSUBS 0.151f
C424 pdrv2.t118 VSUBS 0.151f
C425 pdrv2.t33 VSUBS 0.151f
C426 pdrv2.t189 VSUBS 0.151f
C427 pdrv2.t138 VSUBS 0.151f
C428 pdrv2.t20 VSUBS 0.151f
C429 pdrv2.t62 VSUBS 0.151f
C430 pdrv2.t162 VSUBS 0.151f
C431 pdrv2.t16 VSUBS 0.151f
C432 pdrv2.t49 VSUBS 0.151f
C433 pdrv2.t145 VSUBS 0.151f
C434 pdrv2.t136 VSUBS 0.151f
C435 pdrv2.t32 VSUBS 0.151f
C436 pdrv2.t66 VSUBS 0.151f
C437 pdrv2.t168 VSUBS 0.151f
C438 pdrv2.t22 VSUBS 0.151f
C439 pdrv2.t11 VSUBS 0.151f
C440 pdrv2.t91 VSUBS 0.151f
C441 pdrv2.t21 VSUBS 0.151f
C442 pdrv2.t102 VSUBS 0.151f
C443 pdrv2.n116 VSUBS 0.273f
C444 pdrv2.n117 VSUBS 0.187f
C445 pdrv2.n118 VSUBS 0.187f
C446 pdrv2.n119 VSUBS 0.187f
C447 pdrv2.n120 VSUBS 0.187f
C448 pdrv2.n121 VSUBS 0.187f
C449 pdrv2.n122 VSUBS 0.187f
C450 pdrv2.n123 VSUBS 0.288f
C451 pdrv2.n124 VSUBS 0.324f
C452 pdrv2.n125 VSUBS 0.271f
C453 pdrv2.n126 VSUBS 0.272f
C454 pdrv2.n127 VSUBS 0.177f
C455 pdrv2.n128 VSUBS 0.177f
C456 pdrv2.n129 VSUBS 0.177f
C457 pdrv2.n130 VSUBS 0.177f
C458 pdrv2.n131 VSUBS 0.177f
C459 pdrv2.n132 VSUBS 0.271f
C460 pdrv2.t87 VSUBS 0.151f
C461 pdrv2.t65 VSUBS 0.151f
C462 pdrv2.t6 VSUBS 0.151f
C463 pdrv2.t180 VSUBS 0.151f
C464 pdrv2.t82 VSUBS 0.151f
C465 pdrv2.t57 VSUBS 0.151f
C466 pdrv2.t199 VSUBS 0.151f
C467 pdrv2.t169 VSUBS 0.151f
C468 pdrv2.t7 VSUBS 0.151f
C469 pdrv2.t181 VSUBS 0.151f
C470 pdrv2.t156 VSUBS 0.151f
C471 pdrv2.t127 VSUBS 0.151f
C472 pdrv2.t56 VSUBS 0.151f
C473 pdrv2.t38 VSUBS 0.151f
C474 pdrv2.t25 VSUBS 0.151f
C475 pdrv2.t198 VSUBS 0.151f
C476 pdrv2.t120 VSUBS 0.151f
C477 pdrv2.t97 VSUBS 0.151f
C478 pdrv2.t128 VSUBS 0.151f
C479 pdrv2.t104 VSUBS 0.151f
C480 pdrv2.t40 VSUBS 0.151f
C481 pdrv2.t24 VSUBS 0.151f
C482 pdrv2.t1 VSUBS 0.151f
C483 pdrv2.t171 VSUBS 0.151f
C484 pdrv2.t152 VSUBS 0.151f
C485 pdrv2.t119 VSUBS 0.151f
C486 pdrv2.t51 VSUBS 0.151f
C487 pdrv2.t34 VSUBS 0.151f
C488 pdrv2.t4 VSUBS 0.151f
C489 pdrv2.t179 VSUBS 0.151f
C490 pdrv2.t125 VSUBS 0.151f
C491 pdrv2.t99 VSUBS 0.151f
C492 pdrv2.t176 VSUBS 0.151f
C493 pdrv2.t149 VSUBS 0.151f
C494 pdrv2.t28 VSUBS 0.151f
C495 pdrv2.t0 VSUBS 0.151f
C496 pdrv2.t108 VSUBS 0.151f
C497 pdrv2.t83 VSUBS 0.151f
C498 pdrv2.t100 VSUBS 0.151f
C499 pdrv2.t76 VSUBS 0.151f
C500 pdrv2.t8 VSUBS 0.151f
C501 pdrv2.t182 VSUBS 0.151f
C502 pdrv2.t52 VSUBS 0.151f
C503 pdrv2.t35 VSUBS 0.151f
C504 pdrv2.t153 VSUBS 0.151f
C505 pdrv2.t122 VSUBS 0.151f
C506 pdrv2.t2 VSUBS 0.151f
C507 pdrv2.t172 VSUBS 0.151f
C508 pdrv2.t194 VSUBS 0.151f
C509 pdrv2.t166 VSUBS 0.151f
C510 pdrv2.t77 VSUBS 0.151f
C511 pdrv2.t54 VSUBS 0.151f
C512 pdrv2.t121 VSUBS 0.151f
C513 pdrv2.t98 VSUBS 0.151f
C514 pdrv2.t84 VSUBS 0.151f
C515 pdrv2.t59 VSUBS 0.151f
C516 pdrv2.t129 VSUBS 0.151f
C517 pdrv2.t103 VSUBS 0.151f
C518 pdrv2.t183 VSUBS 0.151f
C519 pdrv2.t155 VSUBS 0.151f
C520 pdrv2.t29 VSUBS 0.151f
C521 pdrv2.t3 VSUBS 0.151f
C522 pdrv2.t60 VSUBS 0.151f
C523 pdrv2.t43 VSUBS 0.151f
C524 pdrv2.t161 VSUBS 0.151f
C525 pdrv2.t131 VSUBS 0.151f
C526 pdrv2.t67 VSUBS 0.151f
C527 pdrv2.t47 VSUBS 0.151f
C528 pdrv2.t111 VSUBS 0.151f
C529 pdrv2.t85 VSUBS 0.151f
C530 pdrv2.t159 VSUBS 0.151f
C531 pdrv2.t130 VSUBS 0.151f
C532 pdrv2.t185 VSUBS 0.151f
C533 pdrv2.t69 VSUBS 0.151f
C534 pdrv2.t114 VSUBS 0.151f
C535 pdrv2.t164 VSUBS 0.151f
C536 pdrv2.n133 VSUBS 0.266f
C537 pdrv2.n134 VSUBS 0.177f
C538 pdrv2.n135 VSUBS 0.177f
C539 pdrv2.n136 VSUBS 0.177f
C540 pdrv2.n137 VSUBS 0.177f
C541 pdrv2.n138 VSUBS 0.177f
C542 pdrv2.n139 VSUBS 0.177f
C543 pdrv2.n140 VSUBS 0.177f
C544 pdrv2.n141 VSUBS 0.177f
C545 pdrv2.n142 VSUBS 0.177f
C546 pdrv2.n143 VSUBS 0.177f
C547 pdrv2.n144 VSUBS 0.177f
C548 pdrv2.n145 VSUBS 0.177f
C549 pdrv2.n146 VSUBS 0.177f
C550 pdrv2.n147 VSUBS 0.177f
C551 pdrv2.n148 VSUBS 0.177f
C552 pdrv2.n149 VSUBS 0.177f
C553 pdrv2.n150 VSUBS 0.177f
C554 pdrv2.n151 VSUBS 0.177f
C555 pdrv2.n152 VSUBS 0.177f
C556 pdrv2.n153 VSUBS 0.177f
C557 pdrv2.n154 VSUBS 0.177f
C558 pdrv2.n155 VSUBS 0.177f
C559 pdrv2.n156 VSUBS 0.177f
C560 pdrv2.n157 VSUBS 0.177f
C561 pdrv2.n158 VSUBS 0.177f
C562 pdrv2.n159 VSUBS 0.177f
C563 pdrv2.n160 VSUBS 0.177f
C564 pdrv2.n161 VSUBS 0.177f
C565 pdrv2.n162 VSUBS 0.177f
C566 pdrv2.n163 VSUBS 0.177f
C567 pdrv2.t12 VSUBS 0.151f
C568 pdrv2.n164 VSUBS 0.177f
C569 pdrv2.t92 VSUBS 0.151f
C570 pdrv2.n165 VSUBS 0.177f
C571 pdrv2.t141 VSUBS 0.151f
C572 pdrv2.n166 VSUBS 0.177f
C573 pdrv2.t192 VSUBS 0.151f
C574 pdrv2.n167 VSUBS 0.189f
C575 pdrv2.n168 VSUBS 1.36f
C576 VSS.n1 VSUBS 0.0148f
C577 VSS.n2 VSUBS 0.0199f
C578 VSS.n3 VSUBS 0.0148f
C579 VSS.n4 VSUBS 0.0199f
C580 VSS.n6 VSUBS 0.0163f
C581 VSS.n7 VSUBS 0.0268f
C582 VSS.n8 VSUBS 0.042f
C583 VSS.n9 VSUBS 0.0402f
C584 VSS.n10 VSUBS 0.0163f
C585 VSS.n11 VSUBS 0.0268f
C586 VSS.n13 VSUBS 0.0148f
C587 VSS.n14 VSUBS 0.0199f
C588 VSS.n15 VSUBS 0.0148f
C589 VSS.n16 VSUBS 0.0199f
C590 VSS.n18 VSUBS 0.0163f
C591 VSS.n19 VSUBS 0.0268f
C592 VSS.n20 VSUBS 0.0236f
C593 VSS.n21 VSUBS 0.0137f
C594 VSS.n22 VSUBS 0.042f
C595 VSS.n23 VSUBS 0.0402f
C596 VSS.n24 VSUBS 0.0163f
C597 VSS.n25 VSUBS 0.0268f
C598 VSS.n27 VSUBS 0.0148f
C599 VSS.n28 VSUBS 0.0199f
C600 VSS.n29 VSUBS 0.0148f
C601 VSS.n30 VSUBS 0.0199f
C602 VSS.n32 VSUBS 1.15f
C603 VSS.n33 VSUBS 20.8f
C604 VSS.n35 VSUBS 0.0326f
C605 VSS.n36 VSUBS 0.0292f
C606 VSS.n37 VSUBS 0.859f
C607 VSS.n38 VSUBS 0.417f
C608 VSS.n39 VSUBS 1.54f
C609 VSS.n41 VSUBS 0.0184f
C610 VSS.n42 VSUBS 0.00625f
C611 VSS.n43 VSUBS 0.7f
C612 VSS.n44 VSUBS 0.603f
C613 VSS.n45 VSUBS 0.0184f
C614 VSS.n46 VSUBS 0.0103f
C615 VSS.n47 VSUBS 0.0876f
C616 VSS.n48 VSUBS 0.0331f
C617 VSS.n49 VSUBS 0.0703f
C618 VSS.n50 VSUBS 0.139f
C619 VSS.n51 VSUBS 0.859f
C620 VSS.n52 VSUBS 0.0148f
C621 VSS.n53 VSUBS 0.0556f
C622 VSS.n54 VSUBS 0.556f
C623 VSS.n55 VSUBS 0.0186f
C624 VSS.n56 VSUBS 0.0478f
C625 VSS.n57 VSUBS 0.0148f
C626 VSS.n58 VSUBS 0.0478f
C627 VSS.n59 VSUBS 0.0186f
C628 VSS.n60 VSUBS 0.0478f
C629 VSS.n61 VSUBS 0.0148f
C630 VSS.n62 VSUBS 0.0591f
C631 VSS.n63 VSUBS 0.0148f
C632 VSS.n64 VSUBS 0.0256f
C633 VSS.t11 VSUBS 0.72f
C634 VSS.n65 VSUBS 0.303f
C635 VSS.n66 VSUBS 0.139f
C636 VSS.n67 VSUBS 0.417f
C637 VSS.t1 VSUBS 0.303f
C638 VSS.t5 VSUBS 0.429f
C639 VSS.n68 VSUBS 0.429f
C640 VSS.n69 VSUBS 0.682f
C641 VSS.n70 VSUBS 0.846f
C642 VSS.n71 VSUBS 0.859f
C643 VSS.n72 VSUBS 0.189f
C644 VSS.n73 VSUBS 0.0148f
C645 VSS.n74 VSUBS 1.55f
C646 VSS.n75 VSUBS 0.859f
C647 VSS.n76 VSUBS 0.0331f
C648 VSS.n78 VSUBS 0.0185f
C649 VSS.n79 VSUBS 0.022f
C650 VSS.n80 VSUBS 0.0115f
C651 VSS.n81 VSUBS 0.0123f
C652 VSS.n82 VSUBS 0.03f
C653 VSS.n84 VSUBS 0.0148f
C654 VSS.n85 VSUBS 0.045f
C655 VSS.n86 VSUBS 0.0335f
C656 VSS.n87 VSUBS 0.015f
C657 VSS.n88 VSUBS 0.0264f
C658 VSS.n89 VSUBS 0.0148f
C659 VSS.n90 VSUBS 0.045f
C660 VSS.n91 VSUBS 0.0353f
C661 VSS.n93 VSUBS 0.0148f
C662 VSS.n94 VSUBS 0.103f
C663 VSS.n95 VSUBS 0.0148f
C664 VSS.n96 VSUBS 0.0758f
C665 VSS.n97 VSUBS 0.0599f
C666 VSS.n99 VSUBS 0.0148f
C667 VSS.n100 VSUBS 0.0635f
C668 VSS.n101 VSUBS 0.0599f
C669 VSS.n103 VSUBS 0.0148f
C670 VSS.n104 VSUBS 0.0617f
C671 VSS.n105 VSUBS 0.0229f
C672 VSS.n106 VSUBS 0.00353f
C673 VSS.n107 VSUBS 0.0203f
C674 VSS.n108 VSUBS 0.456f
C675 VSS.n109 VSUBS 0.0184f
C676 VSS.n110 VSUBS 0.0599f
C677 VSS.n111 VSUBS 0.0148f
C678 VSS.n112 VSUBS 0.0599f
C679 VSS.n114 VSUBS 0.0184f
C680 VSS.n115 VSUBS 0.0599f
C681 VSS.n116 VSUBS 0.0148f
C682 VSS.n117 VSUBS 0.0767f
C683 VSS.n119 VSUBS 0.0148f
C684 VSS.n120 VSUBS 0.12f
C685 VSS.n121 VSUBS 0.0148f
C686 VSS.n122 VSUBS 0.112f
C687 VSS.n123 VSUBS 0.0186f
C688 VSS.n124 VSUBS 0.124f
C689 VSS.n125 VSUBS 0.0389f
C690 VSS.n126 VSUBS 0.0186f
C691 VSS.n127 VSUBS 0.0586f
C692 VSS.n128 VSUBS 0.0148f
C693 VSS.n129 VSUBS 0.0115f
C694 VSS.n130 VSUBS 0.0148f
C695 VSS.n131 VSUBS 0.00842f
C696 VSS.n132 VSUBS 0.0148f
C697 VSS.n133 VSUBS 0.00842f
C698 VSS.n134 VSUBS 0.0148f
C699 VSS.n135 VSUBS 0.00842f
C700 VSS.n136 VSUBS 0.0148f
C701 VSS.n137 VSUBS 0.00842f
C702 VSS.n138 VSUBS 0.0148f
C703 VSS.n139 VSUBS 0.00842f
C704 VSS.n140 VSUBS 0.0148f
C705 VSS.n141 VSUBS 0.00842f
C706 VSS.n142 VSUBS 0.0148f
C707 VSS.n143 VSUBS 0.00842f
C708 VSS.n144 VSUBS 0.0148f
C709 VSS.n145 VSUBS 0.00842f
C710 VSS.n146 VSUBS 0.0293f
C711 VSS.n147 VSUBS 0.00928f
C712 VSS.n148 VSUBS 0.0255f
C713 VSS.n149 VSUBS 0.106f
C714 VSS.n151 VSUBS 0.0283f
C715 VSS.n152 VSUBS 0.0934f
C716 VSS.n153 VSUBS 0.0509f
C717 VSS.n154 VSUBS 0.0529f
C718 VSS.n155 VSUBS 1.24f
C719 VSS.t6 VSUBS 0.0109f
C720 VSS.n156 VSUBS 0.0351f
C721 VSS.n157 VSUBS 0.00642f
C722 VSS.n158 VSUBS 0.0073f
C723 VSS.n159 VSUBS 0.0172f
C724 VSS.n160 VSUBS 0.00246f
C725 VSS.n161 VSUBS 0.00439f
C726 VSS.n162 VSUBS 0.00108f
C727 VSS.n163 VSUBS 0.00138f
C728 VSS.n164 VSUBS 0.00923f
C729 VSS.n165 VSUBS 0.0303f
C730 VSS.n166 VSUBS 0.0362f
C731 VSS.n167 VSUBS 0.00424f
C732 VSS.n168 VSUBS 0.0537f
C733 VSS.t9 VSUBS 0.0109f
C734 VSS.t7 VSUBS 0.0109f
C735 VSS.n169 VSUBS 0.0241f
C736 VSS.n170 VSUBS 0.0065f
C737 VSS.n171 VSUBS 0.0073f
C738 VSS.n172 VSUBS 0.0169f
C739 VSS.n173 VSUBS 0.00246f
C740 VSS.n174 VSUBS 0.00443f
C741 VSS.n175 VSUBS 0.00108f
C742 VSS.n176 VSUBS 0.00108f
C743 VSS.n177 VSUBS 0.00939f
C744 VSS.n178 VSUBS 0.0314f
C745 VSS.n179 VSUBS 0.0379f
C746 VSS.n180 VSUBS 0.00408f
C747 VSS.n181 VSUBS 0.054f
C748 VSS.t12 VSUBS 0.0109f
C749 VSS.n182 VSUBS 0.0349f
C750 VSS.n183 VSUBS 0.00659f
C751 VSS.n184 VSUBS 0.0073f
C752 VSS.n185 VSUBS 0.0164f
C753 VSS.n186 VSUBS 0.00246f
C754 VSS.n187 VSUBS 0.00447f
C755 VSS.n188 VSUBS 0.00108f
C756 VSS.n189 VSUBS 9.23e-19
C757 VSS.n190 VSUBS 0.00953f
C758 VSS.n191 VSUBS 0.0322f
C759 VSS.n192 VSUBS 0.0377f
C760 VSS.n193 VSUBS 0.00391f
C761 VSS.n194 VSUBS 0.0542f
C762 VSS.t138 VSUBS 0.0109f
C763 VSS.n195 VSUBS 0.0349f
C764 VSS.n196 VSUBS 0.0066f
C765 VSS.n197 VSUBS 0.0073f
C766 VSS.n198 VSUBS 0.0161f
C767 VSS.n199 VSUBS 0.00246f
C768 VSS.n200 VSUBS 0.00447f
C769 VSS.n201 VSUBS 0.00108f
C770 VSS.n202 VSUBS 7.69e-19
C771 VSS.n203 VSUBS 0.00955f
C772 VSS.n204 VSUBS 0.0326f
C773 VSS.n205 VSUBS 0.037f
C774 VSS.n206 VSUBS 0.00392f
C775 VSS.n207 VSUBS 0.0545f
C776 VSS.n208 VSUBS 0.00992f
C777 VSS.n209 VSUBS 0.00411f
C778 VSS.n210 VSUBS 0.024f
C779 VSS.n211 VSUBS 0.014f
C780 VSS.n212 VSUBS 0.0171f
C781 VSS.n213 VSUBS 0.011f
C782 VSS.n214 VSUBS 0.0171f
C783 VSS.n215 VSUBS 0.011f
C784 VSS.n216 VSUBS 0.0171f
C785 VSS.n217 VSUBS 0.011f
C786 VSS.n218 VSUBS 0.0171f
C787 VSS.n219 VSUBS 0.011f
C788 VSS.n220 VSUBS 0.024f
C789 VSS.n221 VSUBS 0.014f
C790 VSS.n222 VSUBS 0.0269f
C791 VSS.n223 VSUBS 0.0148f
C792 VSS.n224 VSUBS 0.0253f
C793 VSS.n225 VSUBS 0.0149f
C794 VSS.n226 VSUBS 0.00845f
C795 VSS.n227 VSUBS 0.00745f
C796 VSS.n228 VSUBS 0.0029f
C797 VSS.n229 VSUBS 0.00629f
C798 VSS.n230 VSUBS 0.00967f
C799 VSS.n231 VSUBS 0.0109f
C800 VSS.n232 VSUBS 0.0148f
C801 VSS.n233 VSUBS 0.0293f
C802 VSS.n235 VSUBS 0.0148f
C803 VSS.n236 VSUBS 0.0283f
C804 VSS.n237 VSUBS 0.0338f
C805 VSS.n238 VSUBS 0.00581f
C806 VSS.n239 VSUBS 0.00556f
C807 VSS.n240 VSUBS 0.0106f
C808 VSS.n241 VSUBS 0.0109f
C809 VSS.n242 VSUBS 0.00581f
C810 VSS.n244 VSUBS 0.0148f
C811 VSS.n245 VSUBS 0.0273f
C812 VSS.n247 VSUBS 0.0406f
C813 VSS.n248 VSUBS 0.0163f
C814 VSS.n249 VSUBS 0.0189f
C815 VSS.n250 VSUBS 0.0214f
C816 VSS.n251 VSUBS 0.00556f
C817 VSS.n252 VSUBS 0.0106f
C818 VSS.n253 VSUBS 0.00992f
C819 VSS.n254 VSUBS 0.00629f
C820 VSS.n255 VSUBS 0.0148f
C821 VSS.n256 VSUBS 0.0179f
C822 VSS.n257 VSUBS 0.0129f
C823 VSS.n258 VSUBS 0.00845f
C824 VSS.n259 VSUBS 0.0148f
C825 VSS.n260 VSUBS 0.0199f
C826 VSS.n261 VSUBS 0.00845f
C827 VSS.n262 VSUBS 0.0029f
C828 VSS.n263 VSUBS 0.00411f
C829 VSS.n264 VSUBS 0.00967f
C830 VSS.n265 VSUBS 0.00895f
C831 VSS.n266 VSUBS 0.00629f
C832 VSS.n268 VSUBS 0.0148f
C833 VSS.n269 VSUBS 0.0179f
C834 VSS.n270 VSUBS 0.0109f
C835 VSS.n271 VSUBS 0.00845f
C836 VSS.n272 VSUBS 0.0148f
C837 VSS.n273 VSUBS 0.0199f
C838 VSS.n274 VSUBS 0.0104f
C839 VSS.n275 VSUBS 0.00484f
C840 VSS.n276 VSUBS 0.00411f
C841 VSS.n277 VSUBS 0.00871f
C842 VSS.n278 VSUBS 0.00798f
C843 VSS.n279 VSUBS 0.00629f
C844 VSS.n281 VSUBS 0.0326f
C845 VSS.n282 VSUBS 0.0199f
C846 VSS.n283 VSUBS 0.0124f
C847 VSS.n284 VSUBS 0.00677f
C848 VSS.n285 VSUBS 0.00339f
C849 VSS.n286 VSUBS 0.00314f
C850 VSS.n287 VSUBS 0.00774f
C851 VSS.n288 VSUBS 0.0109f
C852 VSS.n289 VSUBS 0.00774f
C853 VSS.n290 VSUBS 0.0372f
C854 VSS.n291 VSUBS 0.00696f
C855 VSS.n292 VSUBS 0.00646f
C856 VSS.n293 VSUBS 0.00695f
C857 VSS.n294 VSUBS 0.0148f
C858 VSS.n295 VSUBS 0.0224f
C859 VSS.n296 VSUBS 0.0248f
C860 VSS.n297 VSUBS 0.00546f
C861 VSS.n299 VSUBS 0.0305f
C862 VSS.n300 VSUBS 0.0269f
C863 VSS.n301 VSUBS 0.0148f
C864 VSS.n302 VSUBS 0.0199f
C865 VSS.n304 VSUBS 0.0148f
C866 VSS.n305 VSUBS 0.0199f
C867 VSS.n307 VSUBS 0.0163f
C868 VSS.n308 VSUBS 0.0268f
C869 VSS.n309 VSUBS 0.0423f
C870 VSS.n310 VSUBS 0.0406f
C871 VSS.n311 VSUBS 0.0163f
C872 VSS.n312 VSUBS 0.0269f
C873 VSS.n314 VSUBS 0.0148f
C874 VSS.n315 VSUBS 0.0199f
C875 VSS.n316 VSUBS 0.0148f
C876 VSS.n317 VSUBS 0.0199f
C877 VSS.n319 VSUBS 0.0326f
C878 VSS.n320 VSUBS 0.0634f
C879 VSS.n321 VSUBS 0.0331f
C880 VSS.n322 VSUBS 0.361f
C881 VSS.n323 VSUBS 0.0148f
C882 VSS.n324 VSUBS 0.136f
C883 VSS.n325 VSUBS 0.0148f
C884 VSS.n326 VSUBS 0.136f
C885 VSS.n327 VSUBS 0.0148f
C886 VSS.n328 VSUBS 0.134f
C887 VSS.n329 VSUBS 0.0148f
C888 VSS.n330 VSUBS 0.135f
C889 VSS.n331 VSUBS 0.0331f
C890 VSS.n332 VSUBS 0.307f
C891 VSS.n333 VSUBS 0.273f
C892 VSS.n334 VSUBS 0.0074f
C893 VSS.n335 VSUBS 0.0148f
C894 VSS.n336 VSUBS 0.0283f
C895 VSS.n337 VSUBS 0.0148f
C896 VSS.n339 VSUBS 0.0148f
C897 VSS.n340 VSUBS 0.00674f
C898 VSS.n341 VSUBS 0.0148f
C899 VSS.n342 VSUBS 0.00689f
C900 VSS.n343 VSUBS 0.0148f
C901 VSS.n344 VSUBS 0.00689f
C902 VSS.n345 VSUBS 0.0148f
C903 VSS.n346 VSUBS 0.00689f
C904 VSS.n347 VSUBS 0.0148f
C905 VSS.n348 VSUBS 0.00689f
C906 VSS.n349 VSUBS 0.0148f
C907 VSS.n350 VSUBS 0.00689f
C908 VSS.n351 VSUBS 0.0148f
C909 VSS.n352 VSUBS 0.00689f
C910 VSS.n353 VSUBS 0.0148f
C911 VSS.n354 VSUBS 0.00689f
C912 VSS.n355 VSUBS 0.0148f
C913 VSS.n356 VSUBS 0.00689f
C914 VSS.n357 VSUBS 0.0293f
C915 VSS.n358 VSUBS 0.00781f
C916 VSS.n359 VSUBS 0.0148f
C917 VSS.n360 VSUBS 0.0074f
C918 VSS.t17 VSUBS 1.72f
C919 VSS.n361 VSUBS 1.72f
C920 VSS.n362 VSUBS 1.72f
C921 VSS.n363 VSUBS 1.72f
C922 VSS.n364 VSUBS 1.72f
C923 VSS.n365 VSUBS 1.72f
C924 VSS.n366 VSUBS 0.985f
C925 VSS.t15 VSUBS 0.859f
C926 VSS.n367 VSUBS 1.59f
C927 VSS.n368 VSUBS 1.72f
C928 VSS.n369 VSUBS 2.11f
C929 VSS.n370 VSUBS 4.15f
C930 VSS.n371 VSUBS 0.0148f
C931 VSS.n372 VSUBS 0.0148f
C932 VSS.n373 VSUBS 0.124f
C933 VSS.n374 VSUBS 0.127f
C934 VSS.n375 VSUBS 0.18f
C935 VSS.n376 VSUBS 0.174f
C936 VSS.n377 VSUBS 0.013f
C937 VSS.n378 VSUBS 0.0133f
C938 VSS.n379 VSUBS 0.0118f
C939 VSS.n380 VSUBS 0.00751f
C940 VSS.n381 VSUBS 0.0144f
C941 VSS.n382 VSUBS 0.0162f
C942 VSS.n383 VSUBS 0.00751f
C943 VSS.n384 VSUBS 0.0156f
C944 VSS.n385 VSUBS 0.015f
C945 VSS.n386 VSUBS 0.00751f
C946 VSS.n387 VSUBS 0.0118f
C947 VSS.n388 VSUBS 0.0127f
C948 VSS.n389 VSUBS 0.00664f
C949 VSS.n390 VSUBS 0.00693f
C950 VSS.n391 VSUBS 0.013f
C951 VSS.n392 VSUBS 0.0127f
C952 VSS.n393 VSUBS 0.00664f
C953 VSS.n394 VSUBS 0.00693f
C954 VSS.n395 VSUBS 0.013f
C955 VSS.n396 VSUBS 0.0116f
C956 VSS.n397 VSUBS 0.00751f
C957 VSS.n398 VSUBS 0.0153f
C958 VSS.n399 VSUBS 0.0153f
C959 VSS.n400 VSUBS 0.00751f
C960 VSS.n401 VSUBS 0.0165f
C961 VSS.n402 VSUBS 0.0142f
C962 VSS.n403 VSUBS 0.00375f
C963 VSS.n404 VSUBS 0.0567f
C964 VSS.n405 VSUBS 0.0104f
C965 VSS.n406 VSUBS 0.013f
C966 VSS.n407 VSUBS 0.00871f
C967 VSS.n408 VSUBS 0.00629f
C968 VSS.n409 VSUBS 0.0163f
C969 VSS.n410 VSUBS 0.0184f
C970 VSS.n411 VSUBS 0.0148f
C971 VSS.n412 VSUBS 0.00795f
C972 VSS.n413 VSUBS 0.0129f
C973 VSS.n414 VSUBS 0.00845f
C974 VSS.n415 VSUBS 0.0209f
C975 VSS.n416 VSUBS 0.00483f
C976 VSS.n417 VSUBS 0.00411f
C977 VSS.n418 VSUBS 0.00895f
C978 VSS.n419 VSUBS 0.00774f
C979 VSS.n420 VSUBS 0.00629f
C980 VSS.n421 VSUBS 0.00646f
C981 VSS.n422 VSUBS 0.0219f
C982 VSS.n423 VSUBS 0.00677f
C983 VSS.n424 VSUBS 0.00314f
C984 VSS.n425 VSUBS 0.00339f
C985 VSS.n426 VSUBS 0.00696f
C986 VSS.n428 VSUBS 0.0148f
C987 VSS.n429 VSUBS 0.0184f
C988 VSS.n431 VSUBS 0.0148f
C989 VSS.n432 VSUBS 0.00497f
C990 VSS.n433 VSUBS 0.00895f
C991 VSS.n434 VSUBS 0.00774f
C992 VSS.n435 VSUBS 0.00339f
C993 VSS.n436 VSUBS 0.00314f
C994 VSS.n437 VSUBS 0.00646f
C995 VSS.n438 VSUBS 0.0219f
C996 VSS.n439 VSUBS 0.00774f
C997 VSS.n440 VSUBS 0.0109f
C998 VSS.n441 VSUBS 0.013f
C999 VSS.n442 VSUBS 0.0133f
C1000 VSS.n443 VSUBS 0.0118f
C1001 VSS.n444 VSUBS 0.00751f
C1002 VSS.n445 VSUBS 0.0144f
C1003 VSS.n446 VSUBS 0.0162f
C1004 VSS.n447 VSUBS 0.00751f
C1005 VSS.n448 VSUBS 0.0156f
C1006 VSS.n449 VSUBS 0.015f
C1007 VSS.n450 VSUBS 0.00751f
C1008 VSS.n451 VSUBS 0.0118f
C1009 VSS.n452 VSUBS 0.0127f
C1010 VSS.n453 VSUBS 0.00664f
C1011 VSS.n454 VSUBS 0.00693f
C1012 VSS.n455 VSUBS 0.013f
C1013 VSS.n456 VSUBS 0.0127f
C1014 VSS.n457 VSUBS 0.00664f
C1015 VSS.n458 VSUBS 0.00693f
C1016 VSS.n459 VSUBS 0.013f
C1017 VSS.n460 VSUBS 0.00895f
C1018 VSS.n461 VSUBS 0.0554f
C1019 VSS.n462 VSUBS 0.00578f
C1020 VSS.n463 VSUBS 0.0153f
C1021 VSS.n464 VSUBS 0.0153f
C1022 VSS.n465 VSUBS 0.00751f
C1023 VSS.n466 VSUBS 0.0165f
C1024 VSS.n467 VSUBS 0.0142f
C1025 VSS.n468 VSUBS 0.00751f
C1026 VSS.n469 VSUBS 0.0121f
C1027 VSS.n470 VSUBS 0.013f
C1028 VSS.n471 VSUBS 0.00696f
C1029 VSS.n472 VSUBS 0.0148f
C1030 VSS.n473 VSUBS 0.0214f
C1031 VSS.n474 VSUBS 0.0148f
C1032 VSS.n475 VSUBS 0.00497f
C1033 VSS.n476 VSUBS 0.00895f
C1034 VSS.n477 VSUBS 0.00677f
C1035 VSS.n478 VSUBS 0.00629f
C1036 VSS.n479 VSUBS 0.00798f
C1037 VSS.n480 VSUBS 0.00871f
C1038 VSS.n481 VSUBS 0.00411f
C1039 VSS.n482 VSUBS 0.0258f
C1040 VSS.n483 VSUBS 0.00845f
C1041 VSS.n485 VSUBS 0.0305f
C1042 VSS.n486 VSUBS 0.0214f
C1043 VSS.n488 VSUBS 0.0148f
C1044 VSS.n489 VSUBS 0.00497f
C1045 VSS.n490 VSUBS 0.00696f
C1046 VSS.n491 VSUBS 0.00484f
C1047 VSS.n492 VSUBS 0.00629f
C1048 VSS.n493 VSUBS 0.00895f
C1049 VSS.n494 VSUBS 0.00967f
C1050 VSS.n495 VSUBS 0.00411f
C1051 VSS.n496 VSUBS 0.0278f
C1052 VSS.n497 VSUBS 0.00845f
C1053 VSS.n499 VSUBS 0.0148f
C1054 VSS.n500 VSUBS 0.0288f
C1055 VSS.n501 VSUBS 0.00497f
C1056 VSS.n502 VSUBS 0.0029f
C1057 VSS.n503 VSUBS 0.00629f
C1058 VSS.n504 VSUBS 0.00992f
C1059 VSS.n505 VSUBS 0.0106f
C1060 VSS.n506 VSUBS 0.0148f
C1061 VSS.n507 VSUBS 0.0201f
C1062 VSS.n508 VSUBS 0.0148f
C1063 VSS.n509 VSUBS 0.0201f
C1064 VSS.n511 VSUBS 0.0148f
C1065 VSS.n512 VSUBS 0.0201f
C1066 VSS.n514 VSUBS 0.0148f
C1067 VSS.n515 VSUBS 0.0201f
C1068 VSS.n516 VSUBS 0.0148f
C1069 VSS.n517 VSUBS 0.0201f
C1070 VSS.n519 VSUBS 0.0303f
C1071 VSS.n520 VSUBS 0.027f
C1072 VSS.n521 VSUBS 0.0425f
C1073 VSS.n522 VSUBS 0.0344f
C1074 VSS.n523 VSUBS 0.014f
C1075 VSS.n524 VSUBS 0.0125f
C1076 VSS.n525 VSUBS 0.011f
C1077 VSS.n526 VSUBS 0.00928f
C1078 VSS.n527 VSUBS 0.011f
C1079 VSS.n528 VSUBS 0.0142f
C1080 VSS.n529 VSUBS 0.0143f
C1081 VSS.n530 VSUBS 0.00937f
C1082 VSS.n531 VSUBS 0.011f
C1083 VSS.n532 VSUBS 0.0125f
C1084 VSS.n533 VSUBS 0.011f
C1085 VSS.n534 VSUBS 0.0342f
C1086 VSS.n535 VSUBS 0.0139f
C1087 VSS.n536 VSUBS 0.0393f
C1088 VSS.n537 VSUBS 0.0148f
C1089 VSS.n538 VSUBS 0.0357f
C1090 VSS.n539 VSUBS 0.00895f
C1091 VSS.n540 VSUBS 0.00556f
C1092 VSS.n541 VSUBS 0.00581f
C1093 VSS.n542 VSUBS 0.0109f
C1094 VSS.n543 VSUBS 0.0106f
C1095 VSS.n544 VSUBS 0.00556f
C1096 VSS.n546 VSUBS 0.0303f
C1097 VSS.n547 VSUBS 0.0337f
C1098 VSS.n549 VSUBS 0.0148f
C1099 VSS.n550 VSUBS 0.0149f
C1100 VSS.n551 VSUBS 0.0337f
C1101 VSS.n552 VSUBS 0.00581f
C1102 VSS.n553 VSUBS 0.0109f
C1103 VSS.n554 VSUBS 0.00967f
C1104 VSS.n555 VSUBS 0.00629f
C1105 VSS.n556 VSUBS 0.0148f
C1106 VSS.n557 VSUBS 0.0203f
C1107 VSS.n558 VSUBS 0.0148f
C1108 VSS.n559 VSUBS 0.0248f
C1109 VSS.n560 VSUBS 0.0129f
C1110 VSS.n561 VSUBS 0.00842f
C1111 VSS.n562 VSUBS 9.9e-19
C1112 VSS.n563 VSUBS 0.0029f
C1113 VSS.n564 VSUBS 0.00411f
C1114 VSS.n565 VSUBS 0.00992f
C1115 VSS.n566 VSUBS 0.00871f
C1116 VSS.n567 VSUBS 0.00629f
C1117 VSS.n569 VSUBS 0.0148f
C1118 VSS.n570 VSUBS 0.0203f
C1119 VSS.n572 VSUBS 0.0148f
C1120 VSS.n573 VSUBS 0.0248f
C1121 VSS.n574 VSUBS 0.0109f
C1122 VSS.n575 VSUBS 0.00842f
C1123 VSS.n576 VSUBS 0.00297f
C1124 VSS.n577 VSUBS 0.00483f
C1125 VSS.n578 VSUBS 0.00411f
C1126 VSS.n579 VSUBS 0.00895f
C1127 VSS.n580 VSUBS 0.00774f
C1128 VSS.n581 VSUBS 0.00629f
C1129 VSS.n582 VSUBS 0.0148f
C1130 VSS.n583 VSUBS 0.0203f
C1131 VSS.n584 VSUBS 0.00644f
C1132 VSS.n585 VSUBS 0.00495f
C1133 VSS.n586 VSUBS 0.00677f
C1134 VSS.n587 VSUBS 0.00314f
C1135 VSS.n588 VSUBS 0.00339f
C1136 VSS.n589 VSUBS 0.00693f
C1137 VSS.n590 VSUBS 0.0148f
C1138 VSS.n591 VSUBS 0.0218f
C1139 VSS.n592 VSUBS 0.00693f
C1140 VSS.n593 VSUBS 0.00774f
C1141 VSS.n594 VSUBS 0.0109f
C1142 VSS.n595 VSUBS 0.013f
C1143 VSS.n596 VSUBS 0.0133f
C1144 VSS.n597 VSUBS 0.0118f
C1145 VSS.n598 VSUBS 0.00751f
C1146 VSS.n599 VSUBS 0.0144f
C1147 VSS.n600 VSUBS 0.0133f
C1148 VSS.n601 VSUBS 0.0549f
C1149 VSS.n602 VSUBS 0.00635f
C1150 VSS.n603 VSUBS 0.0156f
C1151 VSS.n604 VSUBS 0.015f
C1152 VSS.n605 VSUBS 0.00751f
C1153 VSS.n606 VSUBS 0.0118f
C1154 VSS.n607 VSUBS 0.0127f
C1155 VSS.n608 VSUBS 0.00664f
C1156 VSS.n609 VSUBS 0.00693f
C1157 VSS.n610 VSUBS 0.013f
C1158 VSS.n611 VSUBS 0.0127f
C1159 VSS.n612 VSUBS 0.00664f
C1160 VSS.n613 VSUBS 0.00693f
C1161 VSS.n614 VSUBS 0.013f
C1162 VSS.n615 VSUBS 0.0116f
C1163 VSS.n616 VSUBS 0.00751f
C1164 VSS.n617 VSUBS 0.0153f
C1165 VSS.n618 VSUBS 0.0127f
C1166 VSS.n619 VSUBS 0.0539f
C1167 VSS.n620 VSUBS 0.00693f
C1168 VSS.n621 VSUBS 0.0165f
C1169 VSS.n622 VSUBS 0.0142f
C1170 VSS.n623 VSUBS 0.00751f
C1171 VSS.n624 VSUBS 0.0121f
C1172 VSS.n625 VSUBS 0.013f
C1173 VSS.n626 VSUBS 0.013f
C1174 VSS.n627 VSUBS 0.0133f
C1175 VSS.n628 VSUBS 0.0118f
C1176 VSS.n629 VSUBS 0.00751f
C1177 VSS.n630 VSUBS 0.0144f
C1178 VSS.n631 VSUBS 0.0162f
C1179 VSS.n632 VSUBS 0.00751f
C1180 VSS.n633 VSUBS 0.0156f
C1181 VSS.n634 VSUBS 0.015f
C1182 VSS.n635 VSUBS 0.00751f
C1183 VSS.n636 VSUBS 0.0118f
C1184 VSS.n637 VSUBS 0.0127f
C1185 VSS.n638 VSUBS 0.00664f
C1186 VSS.n639 VSUBS 0.00693f
C1187 VSS.n640 VSUBS 0.013f
C1188 VSS.n641 VSUBS 0.0127f
C1189 VSS.n642 VSUBS 0.00664f
C1190 VSS.n643 VSUBS 0.00693f
C1191 VSS.n644 VSUBS 0.0158f
C1192 VSS.n645 VSUBS 0.00872f
C1193 VSS.n646 VSUBS 0.0203f
C1194 VSS.n647 VSUBS 0.00767f
C1195 VSS.n648 VSUBS 0.0176f
C1196 VSS.n649 VSUBS 0.0165f
C1197 VSS.n650 VSUBS 0.0142f
C1198 VSS.n651 VSUBS 0.00751f
C1199 VSS.n652 VSUBS 0.0121f
C1200 VSS.n653 VSUBS 0.013f
C1201 VSS.t4 VSUBS 0.0228f
C1202 VSS.t3 VSUBS 0.0229f
C1203 VSS.n654 VSUBS 0.412f
C1204 VSS.n655 VSUBS 0.0863f
C1205 VSS.n656 VSUBS 0.0299f
C1206 VSS.n657 VSUBS 0.0248f
C1207 VSS.n658 VSUBS 0.0148f
C1208 VSS.n659 VSUBS 0.0199f
C1209 VSS.n661 VSUBS 0.0402f
C1210 VSS.n662 VSUBS 0.0163f
C1211 VSS.n663 VSUBS 0.0268f
C1212 VSS.n664 VSUBS 0.0148f
C1213 VSS.n665 VSUBS 0.0199f
C1214 VSS.n667 VSUBS 0.0163f
C1215 VSS.n668 VSUBS 0.0268f
C1216 VSS.n669 VSUBS 0.042f
C1217 VSS.n670 VSUBS 0.0236f
C1218 VSS.n671 VSUBS 0.0137f
C1219 VSS.n672 VSUBS 0.0168f
C1220 VSS.n673 VSUBS 0.0107f
C1221 VSS.n674 VSUBS 0.0168f
C1222 VSS.n675 VSUBS 0.0107f
C1223 VSS.n676 VSUBS 0.0168f
C1224 VSS.n677 VSUBS 0.0107f
C1225 VSS.n678 VSUBS 0.0168f
C1226 VSS.n679 VSUBS 0.0107f
C1227 VSS.n680 VSUBS 0.0236f
C1228 VSS.n681 VSUBS 0.0137f
C1229 VSS.n682 VSUBS 0.0337f
C1230 VSS.n683 VSUBS 0.0154f
C1231 VSS.n685 VSUBS 0.0148f
C1232 VSS.n686 VSUBS 0.00833f
C1233 VSS.n687 VSUBS 0.0337f
C1234 VSS.n688 VSUBS 0.0148f
C1235 VSS.n689 VSUBS 0.00766f
C1236 VSS.n690 VSUBS 0.0184f
C1237 VSS.n691 VSUBS 0.00658f
C1238 VSS.n693 VSUBS 0.0148f
C1239 VSS.n694 VSUBS 0.0203f
C1240 VSS.n695 VSUBS 0.00644f
C1241 VSS.n696 VSUBS 0.00495f
C1242 VSS.n697 VSUBS 0.00774f
C1243 VSS.n698 VSUBS 0.00314f
C1244 VSS.n699 VSUBS 0.00339f
C1245 VSS.n700 VSUBS 0.00693f
C1246 VSS.n702 VSUBS 0.0148f
C1247 VSS.n703 VSUBS 0.0218f
C1248 VSS.n704 VSUBS 0.00693f
C1249 VSS.n705 VSUBS 0.00677f
C1250 VSS.n706 VSUBS 0.00629f
C1251 VSS.n707 VSUBS 0.00798f
C1252 VSS.n708 VSUBS 0.00871f
C1253 VSS.n709 VSUBS 0.00411f
C1254 VSS.n710 VSUBS 0.0148f
C1255 VSS.n711 VSUBS 0.0233f
C1256 VSS.n712 VSUBS 0.00891f
C1257 VSS.n713 VSUBS 0.00842f
C1258 VSS.n714 VSUBS 0.0148f
C1259 VSS.n715 VSUBS 0.0218f
C1260 VSS.n716 VSUBS 0.00495f
C1261 VSS.n717 VSUBS 0.00484f
C1262 VSS.n718 VSUBS 0.00629f
C1263 VSS.n719 VSUBS 0.00895f
C1264 VSS.n720 VSUBS 0.00967f
C1265 VSS.n721 VSUBS 0.00411f
C1266 VSS.n723 VSUBS 0.0148f
C1267 VSS.n724 VSUBS 0.0233f
C1268 VSS.n725 VSUBS 0.0109f
C1269 VSS.n726 VSUBS 0.00842f
C1270 VSS.n728 VSUBS 0.0148f
C1271 VSS.n729 VSUBS 0.0218f
C1272 VSS.n730 VSUBS 0.00297f
C1273 VSS.n731 VSUBS 0.0029f
C1274 VSS.n732 VSUBS 0.00629f
C1275 VSS.n733 VSUBS 0.00992f
C1276 VSS.n734 VSUBS 0.0106f
C1277 VSS.n736 VSUBS 0.0148f
C1278 VSS.n737 VSUBS 0.0327f
C1279 VSS.n738 VSUBS 0.0148f
C1280 VSS.n739 VSUBS 0.0208f
C1281 VSS.n740 VSUBS 0.0139f
C1282 VSS.n741 VSUBS 0.00556f
C1283 VSS.n742 VSUBS 0.00581f
C1284 VSS.n743 VSUBS 0.0109f
C1285 VSS.n744 VSUBS 0.0106f
C1286 VSS.n745 VSUBS 0.00556f
C1287 VSS.n746 VSUBS 0.0148f
C1288 VSS.n747 VSUBS 0.0337f
C1289 VSS.n749 VSUBS 0.0148f
C1290 VSS.n750 VSUBS 0.0149f
C1291 VSS.n752 VSUBS 0.0148f
C1292 VSS.n753 VSUBS 0.0327f
C1293 VSS.n754 VSUBS 0.0198f
C1294 VSS.n755 VSUBS 0.00581f
C1295 VSS.n756 VSUBS 0.0109f
C1296 VSS.n757 VSUBS 0.00967f
C1297 VSS.n758 VSUBS 0.00629f
C1298 VSS.n759 VSUBS 0.0148f
C1299 VSS.n760 VSUBS 0.0163f
C1300 VSS.n761 VSUBS 0.0168f
C1301 VSS.n762 VSUBS 0.00842f
C1302 VSS.n763 VSUBS 0.00297f
C1303 VSS.n764 VSUBS 0.0029f
C1304 VSS.n765 VSUBS 0.00411f
C1305 VSS.n766 VSUBS 0.00992f
C1306 VSS.n767 VSUBS 0.00871f
C1307 VSS.n768 VSUBS 0.00629f
C1308 VSS.n769 VSUBS 0.0148f
C1309 VSS.n770 VSUBS 0.0228f
C1310 VSS.n772 VSUBS 0.0292f
C1311 VSS.n773 VSUBS 0.0163f
C1312 VSS.n774 VSUBS 0.0149f
C1313 VSS.n775 VSUBS 0.00842f
C1314 VSS.n776 VSUBS 0.00495f
C1315 VSS.n777 VSUBS 0.00483f
C1316 VSS.n778 VSUBS 0.00411f
C1317 VSS.n779 VSUBS 0.00895f
C1318 VSS.n780 VSUBS 0.00774f
C1319 VSS.n781 VSUBS 0.00629f
C1320 VSS.n783 VSUBS 0.0148f
C1321 VSS.n784 VSUBS 0.0252f
C1322 VSS.n785 VSUBS 0.00644f
C1323 VSS.n786 VSUBS 0.0208f
C1324 VSS.n787 VSUBS 0.00677f
C1325 VSS.n788 VSUBS 0.00314f
C1326 VSS.n789 VSUBS 0.00339f
C1327 VSS.n790 VSUBS 0.00693f
C1328 VSS.n791 VSUBS 0.0148f
C1329 VSS.n792 VSUBS 0.0201f
C1330 VSS.n793 VSUBS 0.0148f
C1331 VSS.n794 VSUBS 0.0201f
C1332 VSS.n796 VSUBS 0.0148f
C1333 VSS.n797 VSUBS 0.0201f
C1334 VSS.n798 VSUBS 0.0148f
C1335 VSS.n799 VSUBS 0.0201f
C1336 VSS.n801 VSUBS 0.0292f
C1337 VSS.n802 VSUBS 0.027f
C1338 VSS.n803 VSUBS 0.0148f
C1339 VSS.n804 VSUBS 0.0199f
C1340 VSS.n806 VSUBS 0.0294f
C1341 VSS.n807 VSUBS 0.0266f
C1342 VSS.n808 VSUBS 0.0418f
C1343 VSS.n809 VSUBS 0.0358f
C1344 VSS.n810 VSUBS 0.0134f
C1345 VSS.n811 VSUBS 0.013f
C1346 VSS.n812 VSUBS 0.0105f
C1347 VSS.n813 VSUBS 0.00966f
C1348 VSS.n814 VSUBS 0.0105f
C1349 VSS.n815 VSUBS 0.0118f
C1350 VSS.n816 VSUBS 0.0119f
C1351 VSS.n817 VSUBS 0.00976f
C1352 VSS.n818 VSUBS 0.0105f
C1353 VSS.n819 VSUBS 0.013f
C1354 VSS.n820 VSUBS 0.0105f
C1355 VSS.n821 VSUBS 0.0356f
C1356 VSS.n822 VSUBS 0.0133f
C1357 VSS.n823 VSUBS 0.0245f
C1358 VSS.n824 VSUBS 0.0148f
C1359 VSS.n825 VSUBS 0.00895f
C1360 VSS.n826 VSUBS 0.0109f
C1361 VSS.n827 VSUBS 0.00774f
C1362 VSS.n828 VSUBS 0.0109f
C1363 VSS.n829 VSUBS 0.00646f
C1364 VSS.n830 VSUBS 0.0179f
C1365 VSS.n831 VSUBS 0.00774f
C1366 VSS.n832 VSUBS 0.00314f
C1367 VSS.n833 VSUBS 0.00339f
C1368 VSS.n834 VSUBS 0.00696f
C1369 VSS.n835 VSUBS 0.0148f
C1370 VSS.n836 VSUBS 0.0253f
C1371 VSS.n837 VSUBS 0.0109f
C1372 VSS.n838 VSUBS 0.00677f
C1373 VSS.n839 VSUBS 0.00629f
C1374 VSS.n840 VSUBS 0.00798f
C1375 VSS.n841 VSUBS 0.00871f
C1376 VSS.n842 VSUBS 0.00411f
C1377 VSS.n843 VSUBS 0.0248f
C1378 VSS.n844 VSUBS 0.00646f
C1379 VSS.n845 VSUBS 0.0294f
C1380 VSS.n846 VSUBS 0.00298f
C1381 VSS.n848 VSUBS 0.0148f
C1382 VSS.n849 VSUBS 0.0253f
C1383 VSS.n850 VSUBS 0.00795f
C1384 VSS.n851 VSUBS 0.00484f
C1385 VSS.n852 VSUBS 0.00629f
C1386 VSS.n853 VSUBS 0.00895f
C1387 VSS.n854 VSUBS 0.00967f
C1388 VSS.n855 VSUBS 0.00411f
C1389 VSS.n856 VSUBS 0.0258f
C1390 VSS.n858 VSUBS 0.0148f
C1391 VSS.n859 VSUBS 0.00745f
C1392 VSS.n860 VSUBS 0.00199f
C1393 VSS.n861 VSUBS 0.0148f
C1394 VSS.n862 VSUBS 0.0318f
C1395 VSS.n863 VSUBS 0.00696f
C1396 VSS.n864 VSUBS 0.0029f
C1397 VSS.n865 VSUBS 0.00629f
C1398 VSS.n866 VSUBS 0.00992f
C1399 VSS.n867 VSUBS 0.0106f
C1400 VSS.n869 VSUBS 0.0148f
C1401 VSS.n870 VSUBS 0.0288f
C1402 VSS.n872 VSUBS 0.0148f
C1403 VSS.n873 VSUBS 0.0308f
C1404 VSS.n874 VSUBS 0.00795f
C1405 VSS.n875 VSUBS 0.00556f
C1406 VSS.n876 VSUBS 0.00581f
C1407 VSS.n877 VSUBS 0.0109f
C1408 VSS.n878 VSUBS 0.0106f
C1409 VSS.n879 VSUBS 0.00556f
C1410 VSS.n880 VSUBS 0.0402f
C1411 VSS.n881 VSUBS 0.0163f
C1412 VSS.n882 VSUBS 0.0308f
C1413 VSS.n883 VSUBS 0.0148f
C1414 VSS.n884 VSUBS 0.0355f
C1415 VSS.n885 VSUBS 0.00795f
C1416 VSS.n886 VSUBS 0.00581f
C1417 VSS.n887 VSUBS 0.00653f
C1418 VSS.n888 VSUBS 0.0116f
C1419 VSS.n889 VSUBS 0.00629f
C1420 VSS.n890 VSUBS 0.00629f
C1421 VSS.n891 VSUBS 0.00497f
C1422 VSS.n893 VSUBS 0.0148f
C1423 VSS.n894 VSUBS 0.00447f
C1424 VSS.n895 VSUBS 0.03f
C1425 VSS.n896 VSUBS 0.00677f
C1426 VSS.n897 VSUBS 0.00314f
C1427 VSS.n898 VSUBS 0.00339f
C1428 VSS.n900 VSUBS 0.0163f
C1429 VSS.n901 VSUBS 0.00696f
C1430 VSS.n902 VSUBS 0.0273f
C1431 VSS.n903 VSUBS 0.00774f
C1432 VSS.n904 VSUBS 0.00339f
C1433 VSS.n905 VSUBS 0.00314f
C1434 VSS.n906 VSUBS 0.00497f
C1435 VSS.n908 VSUBS 0.0148f
C1436 VSS.n909 VSUBS 0.00447f
C1437 VSS.n910 VSUBS 0.0239f
C1438 VSS.n911 VSUBS 0.00774f
C1439 VSS.n912 VSUBS 0.0109f
C1440 VSS.n913 VSUBS 0.013f
C1441 VSS.n914 VSUBS 0.0133f
C1442 VSS.n915 VSUBS 0.0118f
C1443 VSS.n916 VSUBS 0.00751f
C1444 VSS.n917 VSUBS 0.0144f
C1445 VSS.n918 VSUBS 0.0162f
C1446 VSS.n919 VSUBS 0.00751f
C1447 VSS.n920 VSUBS 0.0156f
C1448 VSS.n921 VSUBS 0.015f
C1449 VSS.n922 VSUBS 0.00751f
C1450 VSS.n923 VSUBS 0.0118f
C1451 VSS.n924 VSUBS 0.0127f
C1452 VSS.n925 VSUBS 0.00664f
C1453 VSS.n926 VSUBS 0.00693f
C1454 VSS.n927 VSUBS 0.013f
C1455 VSS.n928 VSUBS 0.0127f
C1456 VSS.n929 VSUBS 0.00664f
C1457 VSS.n930 VSUBS 0.00693f
C1458 VSS.n931 VSUBS 0.013f
C1459 VSS.n932 VSUBS 0.0116f
C1460 VSS.n933 VSUBS 0.00751f
C1461 VSS.n934 VSUBS 0.0153f
C1462 VSS.n935 VSUBS 0.0153f
C1463 VSS.n936 VSUBS 0.00751f
C1464 VSS.n937 VSUBS 0.0165f
C1465 VSS.n938 VSUBS 0.0142f
C1466 VSS.n939 VSUBS 0.00751f
C1467 VSS.n940 VSUBS 0.0121f
C1468 VSS.n941 VSUBS 0.013f
C1469 VSS.n942 VSUBS 0.0148f
C1470 VSS.n943 VSUBS 0.00696f
C1471 VSS.n944 VSUBS 0.0288f
C1472 VSS.n945 VSUBS 0.00677f
C1473 VSS.n946 VSUBS 0.00629f
C1474 VSS.n947 VSUBS 0.00798f
C1475 VSS.n948 VSUBS 0.00871f
C1476 VSS.n949 VSUBS 0.00411f
C1477 VSS.n950 VSUBS 0.0148f
C1478 VSS.n951 VSUBS 0.0253f
C1479 VSS.n952 VSUBS 0.00497f
C1480 VSS.n953 VSUBS 0.0148f
C1481 VSS.n954 VSUBS 0.00546f
C1482 VSS.n955 VSUBS 0.00497f
C1483 VSS.n956 VSUBS 0.0268f
C1484 VSS.n957 VSUBS 0.00484f
C1485 VSS.n958 VSUBS 0.00629f
C1486 VSS.n959 VSUBS 0.00895f
C1487 VSS.n960 VSUBS 0.00967f
C1488 VSS.n961 VSUBS 0.00411f
C1489 VSS.n962 VSUBS 0.0148f
C1490 VSS.n963 VSUBS 0.0253f
C1491 VSS.n964 VSUBS 0.00497f
C1492 VSS.n966 VSUBS 0.0163f
C1493 VSS.n967 VSUBS 0.00745f
C1494 VSS.n968 VSUBS 0.00497f
C1495 VSS.n969 VSUBS 0.0248f
C1496 VSS.n970 VSUBS 0.0029f
C1497 VSS.n971 VSUBS 0.00629f
C1498 VSS.n972 VSUBS 0.00992f
C1499 VSS.n973 VSUBS 0.0106f
C1500 VSS.n975 VSUBS 0.0148f
C1501 VSS.n976 VSUBS 0.0348f
C1502 VSS.n977 VSUBS 0.0148f
C1503 VSS.n978 VSUBS 0.0199f
C1504 VSS.n980 VSUBS 0.0402f
C1505 VSS.n981 VSUBS 0.0163f
C1506 VSS.n982 VSUBS 0.0268f
C1507 VSS.n983 VSUBS 0.0148f
C1508 VSS.n984 VSUBS 0.0199f
C1509 VSS.n986 VSUBS 0.0163f
C1510 VSS.n987 VSUBS 0.0268f
C1511 VSS.n988 VSUBS 0.042f
C1512 VSS.n989 VSUBS 0.0236f
C1513 VSS.n990 VSUBS 0.0137f
C1514 VSS.n991 VSUBS 0.0168f
C1515 VSS.n992 VSUBS 0.0107f
C1516 VSS.n993 VSUBS 0.0168f
C1517 VSS.n994 VSUBS 0.0107f
C1518 VSS.n995 VSUBS 0.0168f
C1519 VSS.n996 VSUBS 0.0107f
C1520 VSS.n997 VSUBS 0.0168f
C1521 VSS.n998 VSUBS 0.0107f
C1522 VSS.n999 VSUBS 0.0236f
C1523 VSS.n1000 VSUBS 0.0137f
C1524 VSS.n1001 VSUBS 0.0312f
C1525 VSS.n1002 VSUBS 0.0283f
C1526 VSS.n1003 VSUBS 0.00556f
C1527 VSS.n1004 VSUBS 0.00581f
C1528 VSS.n1005 VSUBS 0.0109f
C1529 VSS.n1006 VSUBS 0.0106f
C1530 VSS.n1007 VSUBS 0.00556f
C1531 VSS.n1009 VSUBS 0.0148f
C1532 VSS.n1010 VSUBS 0.0184f
C1533 VSS.n1011 VSUBS 0.0148f
C1534 VSS.n1012 VSUBS 0.0353f
C1535 VSS.n1013 VSUBS 0.0338f
C1536 VSS.n1014 VSUBS 0.00581f
C1537 VSS.n1015 VSUBS 0.0109f
C1538 VSS.n1016 VSUBS 0.00967f
C1539 VSS.n1017 VSUBS 0.00629f
C1540 VSS.n1018 VSUBS 0.0159f
C1541 VSS.n1019 VSUBS 0.0402f
C1542 VSS.n1020 VSUBS 0.0163f
C1543 VSS.n1021 VSUBS 0.00795f
C1544 VSS.n1022 VSUBS 0.00348f
C1545 VSS.n1023 VSUBS 0.0149f
C1546 VSS.n1024 VSUBS 0.0029f
C1547 VSS.n1025 VSUBS 0.00411f
C1548 VSS.n1026 VSUBS 0.00992f
C1549 VSS.n1027 VSUBS 0.00871f
C1550 VSS.n1028 VSUBS 0.00629f
C1551 VSS.n1029 VSUBS 0.0148f
C1552 VSS.n1030 VSUBS 0.0253f
C1553 VSS.n1031 VSUBS 0.0159f
C1554 VSS.n1033 VSUBS 0.0148f
C1555 VSS.n1034 VSUBS 0.00596f
C1556 VSS.n1035 VSUBS 0.00348f
C1557 VSS.n1036 VSUBS 0.0169f
C1558 VSS.n1037 VSUBS 0.00483f
C1559 VSS.n1038 VSUBS 0.00411f
C1560 VSS.n1039 VSUBS 0.00895f
C1561 VSS.n1040 VSUBS 0.00774f
C1562 VSS.n1041 VSUBS 0.00629f
C1563 VSS.n1043 VSUBS 0.0148f
C1564 VSS.n1044 VSUBS 0.0253f
C1565 VSS.n1045 VSUBS 0.00298f
C1566 VSS.n1046 VSUBS 0.0148f
C1567 VSS.n1047 VSUBS 0.00447f
C1568 VSS.n1048 VSUBS 0.0179f
C1569 VSS.n1049 VSUBS 0.00677f
C1570 VSS.n1050 VSUBS 0.00314f
C1571 VSS.n1051 VSUBS 0.00339f
C1572 VSS.n1052 VSUBS 0.00696f
C1573 VSS.n1054 VSUBS 0.0148f
C1574 VSS.n1055 VSUBS 0.0224f
C1575 VSS.n1056 VSUBS 0.0129f
C1576 VSS.n1057 VSUBS 0.00774f
C1577 VSS.n1058 VSUBS 0.00339f
C1578 VSS.n1059 VSUBS 0.00314f
C1579 VSS.n1060 VSUBS 0.00298f
C1580 VSS.n1062 VSUBS 0.0163f
C1581 VSS.n1063 VSUBS 0.00447f
C1582 VSS.n1064 VSUBS 0.0179f
C1583 VSS.n1065 VSUBS 0.00774f
C1584 VSS.n1066 VSUBS 0.0109f
C1585 VSS.n1067 VSUBS 0.013f
C1586 VSS.n1068 VSUBS 0.0133f
C1587 VSS.n1069 VSUBS 0.0118f
C1588 VSS.n1070 VSUBS 0.00751f
C1589 VSS.n1071 VSUBS 0.0144f
C1590 VSS.n1072 VSUBS 0.0162f
C1591 VSS.n1073 VSUBS 0.00751f
C1592 VSS.n1074 VSUBS 0.0156f
C1593 VSS.n1075 VSUBS 0.015f
C1594 VSS.n1076 VSUBS 0.00751f
C1595 VSS.n1077 VSUBS 0.0118f
C1596 VSS.n1078 VSUBS 0.0127f
C1597 VSS.n1079 VSUBS 0.00664f
C1598 VSS.n1080 VSUBS 0.00693f
C1599 VSS.n1081 VSUBS 0.013f
C1600 VSS.n1082 VSUBS 0.0127f
C1601 VSS.n1083 VSUBS 0.00664f
C1602 VSS.n1084 VSUBS 0.00693f
C1603 VSS.n1085 VSUBS 0.013f
C1604 VSS.n1086 VSUBS 0.0116f
C1605 VSS.n1087 VSUBS 0.00751f
C1606 VSS.n1088 VSUBS 0.0153f
C1607 VSS.n1089 VSUBS 0.0153f
C1608 VSS.n1090 VSUBS 0.00751f
C1609 VSS.n1091 VSUBS 0.0165f
C1610 VSS.n1092 VSUBS 0.0142f
C1611 VSS.n1093 VSUBS 0.00751f
C1612 VSS.n1094 VSUBS 0.0121f
C1613 VSS.n1095 VSUBS 0.013f
C1614 VSS.t13 VSUBS 0.0256f
C1615 VSS.n1096 VSUBS 0.00696f
C1616 VSS.n1097 VSUBS 0.0148f
C1617 VSS.n1098 VSUBS 0.0253f
C1618 VSS.n1099 VSUBS 0.0129f
C1619 VSS.n1100 VSUBS 0.00435f
C1620 VSS.n1101 VSUBS 0.233f
C1621 VSS.n1102 VSUBS 0.00435f
C1622 VSS.n1103 VSUBS 0.00798f
C1623 VSS.n1104 VSUBS 0.00871f
C1624 VSS.n1105 VSUBS 0.00411f
C1625 VSS.n1106 VSUBS 0.0229f
C1626 VSS.n1107 VSUBS 0.00845f
C1627 VSS.n1108 VSUBS 0.0148f
C1628 VSS.n1109 VSUBS 0.0199f
C1629 VSS.n1111 VSUBS 0.0163f
C1630 VSS.n1112 VSUBS 0.0268f
C1631 VSS.n1113 VSUBS 0.0148f
C1632 VSS.n1114 VSUBS 0.0199f
C1633 VSS.n1115 VSUBS 0.0402f
C1634 VSS.n1117 VSUBS 0.0163f
C1635 VSS.n1118 VSUBS 0.0268f
C1636 VSS.n1119 VSUBS 0.042f
C1637 VSS.n1120 VSUBS 0.0236f
C1638 VSS.n1121 VSUBS 0.0137f
C1639 VSS.n1122 VSUBS 0.0168f
C1640 VSS.n1123 VSUBS 0.0107f
C1641 VSS.n1124 VSUBS 0.0168f
C1642 VSS.n1125 VSUBS 0.0107f
C1643 VSS.n1126 VSUBS 0.0168f
C1644 VSS.n1127 VSUBS 0.0107f
C1645 VSS.n1128 VSUBS 0.0168f
C1646 VSS.n1129 VSUBS 0.0107f
C1647 VSS.n1130 VSUBS 0.0236f
C1648 VSS.n1131 VSUBS 0.0137f
C1649 VSS.n1132 VSUBS 0.0257f
C1650 VSS.n1133 VSUBS 0.0148f
C1651 VSS.n1134 VSUBS 0.0154f
C1652 VSS.n1135 VSUBS 0.0109f
C1653 VSS.n1136 VSUBS 0.00484f
C1654 VSS.n1137 VSUBS 0.00629f
C1655 VSS.n1138 VSUBS 0.00895f
C1656 VSS.n1139 VSUBS 0.00967f
C1657 VSS.n1140 VSUBS 0.00411f
C1658 VSS.n1141 VSUBS 0.0174f
C1659 VSS.n1142 VSUBS 0.00845f
C1660 VSS.n1144 VSUBS 0.0148f
C1661 VSS.n1145 VSUBS 0.0348f
C1662 VSS.n1146 VSUBS 0.00895f
C1663 VSS.n1147 VSUBS 0.0029f
C1664 VSS.n1148 VSUBS 0.00629f
C1665 VSS.n1149 VSUBS 0.00992f
C1666 VSS.n1150 VSUBS 0.0106f
C1667 VSS.n1151 VSUBS 0.0148f
C1668 VSS.n1152 VSUBS 0.0318f
C1669 VSS.n1153 VSUBS 0.0402f
C1670 VSS.n1154 VSUBS 0.0163f
C1671 VSS.n1155 VSUBS 0.00696f
C1672 VSS.n1156 VSUBS 0.0308f
C1673 VSS.n1157 VSUBS 0.00556f
C1674 VSS.n1158 VSUBS 0.00581f
C1675 VSS.n1159 VSUBS 0.0109f
C1676 VSS.n1160 VSUBS 0.0106f
C1677 VSS.n1161 VSUBS 0.00556f
C1678 VSS.n1163 VSUBS 0.0148f
C1679 VSS.n1164 VSUBS 0.0333f
C1680 VSS.n1166 VSUBS 0.0148f
C1681 VSS.n1167 VSUBS 0.00497f
C1682 VSS.n1168 VSUBS 0.0308f
C1683 VSS.n1169 VSUBS 0.00581f
C1684 VSS.n1170 VSUBS 0.0109f
C1685 VSS.n1171 VSUBS 0.00967f
C1686 VSS.n1172 VSUBS 0.00629f
C1687 VSS.n1173 VSUBS 0.0303f
C1688 VSS.n1174 VSUBS 0.0148f
C1689 VSS.n1175 VSUBS 0.00795f
C1690 VSS.n1176 VSUBS 0.0148f
C1691 VSS.n1177 VSUBS 0.00348f
C1692 VSS.n1178 VSUBS 0.0308f
C1693 VSS.n1179 VSUBS 0.0029f
C1694 VSS.n1180 VSUBS 0.00411f
C1695 VSS.n1181 VSUBS 0.00992f
C1696 VSS.n1182 VSUBS 0.00871f
C1697 VSS.n1183 VSUBS 0.00629f
C1698 VSS.n1184 VSUBS 0.0303f
C1699 VSS.n1186 VSUBS 0.0148f
C1700 VSS.n1187 VSUBS 0.00596f
C1701 VSS.n1188 VSUBS 0.00298f
C1702 VSS.n1190 VSUBS 0.0402f
C1703 VSS.n1191 VSUBS 0.0163f
C1704 VSS.n1192 VSUBS 0.00248f
C1705 VSS.n1193 VSUBS 0.0258f
C1706 VSS.n1194 VSUBS 0.00483f
C1707 VSS.n1195 VSUBS 0.00411f
C1708 VSS.n1196 VSUBS 0.00895f
C1709 VSS.n1197 VSUBS 0.00774f
C1710 VSS.n1198 VSUBS 0.00629f
C1711 VSS.n1199 VSUBS 0.00298f
C1712 VSS.n1200 VSUBS 0.0148f
C1713 VSS.n1201 VSUBS 0.00447f
C1714 VSS.n1202 VSUBS 0.0288f
C1715 VSS.n1203 VSUBS 0.00677f
C1716 VSS.n1204 VSUBS 0.00314f
C1717 VSS.n1205 VSUBS 0.00339f
C1718 VSS.n1206 VSUBS 0.00696f
C1719 VSS.n1207 VSUBS 0.0174f
C1720 VSS.n1208 VSUBS 0.00774f
C1721 VSS.n1209 VSUBS 0.00339f
C1722 VSS.n1210 VSUBS 0.00314f
C1723 VSS.n1211 VSUBS 0.0148f
C1724 VSS.n1212 VSUBS 0.0199f
C1725 VSS.n1214 VSUBS 0.0402f
C1726 VSS.n1215 VSUBS 0.0163f
C1727 VSS.n1216 VSUBS 0.0268f
C1728 VSS.n1217 VSUBS 0.0148f
C1729 VSS.n1218 VSUBS 0.0199f
C1730 VSS.n1220 VSUBS 0.0163f
C1731 VSS.n1221 VSUBS 0.0268f
C1732 VSS.n1222 VSUBS 0.042f
C1733 VSS.n1223 VSUBS 0.0236f
C1734 VSS.n1224 VSUBS 0.0137f
C1735 VSS.n1225 VSUBS 0.0168f
C1736 VSS.n1226 VSUBS 0.0107f
C1737 VSS.n1227 VSUBS 0.0168f
C1738 VSS.n1228 VSUBS 0.0107f
C1739 VSS.n1229 VSUBS 0.0168f
C1740 VSS.n1230 VSUBS 0.0107f
C1741 VSS.n1231 VSUBS 0.0168f
C1742 VSS.n1232 VSUBS 0.0107f
C1743 VSS.n1233 VSUBS 0.0236f
C1744 VSS.n1234 VSUBS 0.0137f
C1745 VSS.n1235 VSUBS 0.0307f
C1746 VSS.n1236 VSUBS 0.00298f
C1747 VSS.n1238 VSUBS 0.0148f
C1748 VSS.n1239 VSUBS 0.00447f
C1749 VSS.n1240 VSUBS 0.0134f
C1750 VSS.n1241 VSUBS 0.00774f
C1751 VSS.n1242 VSUBS 0.0109f
C1752 VSS.n1243 VSUBS 0.013f
C1753 VSS.n1244 VSUBS 0.0133f
C1754 VSS.n1245 VSUBS 0.0118f
C1755 VSS.n1246 VSUBS 0.00751f
C1756 VSS.n1247 VSUBS 0.0144f
C1757 VSS.n1248 VSUBS 0.0162f
C1758 VSS.n1249 VSUBS 0.00751f
C1759 VSS.n1250 VSUBS 0.0156f
C1760 VSS.n1251 VSUBS 0.015f
C1761 VSS.n1252 VSUBS 0.00751f
C1762 VSS.n1253 VSUBS 0.0118f
C1763 VSS.n1254 VSUBS 0.0127f
C1764 VSS.n1255 VSUBS 0.00664f
C1765 VSS.n1256 VSUBS 0.00693f
C1766 VSS.n1257 VSUBS 0.013f
C1767 VSS.n1258 VSUBS 0.0127f
C1768 VSS.n1259 VSUBS 0.00664f
C1769 VSS.n1260 VSUBS 0.00693f
C1770 VSS.n1261 VSUBS 0.013f
C1771 VSS.n1262 VSUBS 0.0116f
C1772 VSS.n1263 VSUBS 0.00751f
C1773 VSS.n1264 VSUBS 0.0153f
C1774 VSS.n1265 VSUBS 0.0153f
C1775 VSS.n1266 VSUBS 0.00751f
C1776 VSS.n1267 VSUBS 0.0165f
C1777 VSS.n1268 VSUBS 0.0142f
C1778 VSS.n1269 VSUBS 0.00751f
C1779 VSS.n1270 VSUBS 0.0121f
C1780 VSS.n1271 VSUBS 0.013f
C1781 VSS.n1272 VSUBS 0.00696f
C1782 VSS.n1273 VSUBS 0.0303f
C1783 VSS.n1274 VSUBS 0.00677f
C1784 VSS.n1275 VSUBS 0.00629f
C1785 VSS.n1276 VSUBS 0.00798f
C1786 VSS.n1277 VSUBS 0.00871f
C1787 VSS.n1278 VSUBS 0.00411f
C1788 VSS.n1279 VSUBS 0.0258f
C1789 VSS.n1280 VSUBS 0.0148f
C1790 VSS.n1281 VSUBS 0.00546f
C1791 VSS.n1282 VSUBS 0.00795f
C1792 VSS.n1283 VSUBS 0.0163f
C1793 VSS.n1284 VSUBS 0.0253f
C1794 VSS.n1285 VSUBS 0.00497f
C1795 VSS.n1286 VSUBS 0.00484f
C1796 VSS.n1287 VSUBS 0.00629f
C1797 VSS.n1288 VSUBS 0.00895f
C1798 VSS.n1289 VSUBS 0.00967f
C1799 VSS.n1290 VSUBS 0.00411f
C1800 VSS.n1291 VSUBS 0.0239f
C1801 VSS.n1293 VSUBS 0.0148f
C1802 VSS.n1294 VSUBS 0.00745f
C1803 VSS.n1295 VSUBS 0.00795f
C1804 VSS.n1297 VSUBS 0.0148f
C1805 VSS.n1298 VSUBS 0.0258f
C1806 VSS.n1299 VSUBS 0.00298f
C1807 VSS.n1300 VSUBS 0.0029f
C1808 VSS.n1301 VSUBS 0.00629f
C1809 VSS.n1302 VSUBS 0.00992f
C1810 VSS.n1303 VSUBS 0.0106f
C1811 VSS.n1305 VSUBS 0.0148f
C1812 VSS.n1306 VSUBS 0.0328f
C1813 VSS.n1307 VSUBS 0.0148f
C1814 VSS.n1308 VSUBS 0.0248f
C1815 VSS.n1309 VSUBS 0.00994f
C1816 VSS.n1310 VSUBS 0.00556f
C1817 VSS.n1311 VSUBS 0.00581f
C1818 VSS.n1312 VSUBS 0.0109f
C1819 VSS.n1313 VSUBS 0.0106f
C1820 VSS.n1314 VSUBS 0.00556f
C1821 VSS.n1315 VSUBS 0.0148f
C1822 VSS.n1316 VSUBS 0.0338f
C1823 VSS.n1318 VSUBS 0.0402f
C1824 VSS.n1319 VSUBS 0.0163f
C1825 VSS.n1320 VSUBS 0.0109f
C1826 VSS.n1322 VSUBS 0.0148f
C1827 VSS.n1323 VSUBS 0.0353f
C1828 VSS.n1324 VSUBS 0.0239f
C1829 VSS.n1325 VSUBS 0.00581f
C1830 VSS.n1326 VSUBS 0.0109f
C1831 VSS.n1327 VSUBS 0.00967f
C1832 VSS.n1328 VSUBS 0.00629f
C1833 VSS.n1329 VSUBS 0.0204f
C1834 VSS.n1330 VSUBS 0.00845f
C1835 VSS.n1331 VSUBS 0.0129f
C1836 VSS.n1332 VSUBS 0.0029f
C1837 VSS.n1333 VSUBS 0.00411f
C1838 VSS.n1334 VSUBS 0.00992f
C1839 VSS.n1335 VSUBS 0.00871f
C1840 VSS.n1336 VSUBS 0.00629f
C1841 VSS.n1337 VSUBS 0.0148f
C1842 VSS.n1338 VSUBS 0.0199f
C1843 VSS.n1340 VSUBS 0.0163f
C1844 VSS.n1341 VSUBS 0.0268f
C1845 VSS.n1342 VSUBS 0.0402f
C1846 VSS.n1343 VSUBS 0.0163f
C1847 VSS.n1344 VSUBS 0.0268f
C1848 VSS.n1345 VSUBS 0.042f
C1849 VSS.n1346 VSUBS 0.0236f
C1850 VSS.n1347 VSUBS 0.0137f
C1851 VSS.n1348 VSUBS 0.0168f
C1852 VSS.n1349 VSUBS 0.0107f
C1853 VSS.n1350 VSUBS 0.0168f
C1854 VSS.n1351 VSUBS 0.0107f
C1855 VSS.n1352 VSUBS 0.0168f
C1856 VSS.n1353 VSUBS 0.0107f
C1857 VSS.n1354 VSUBS 0.0168f
C1858 VSS.n1355 VSUBS 0.0107f
C1859 VSS.n1356 VSUBS 0.0236f
C1860 VSS.n1357 VSUBS 0.0137f
C1861 VSS.n1358 VSUBS 0.0213f
C1862 VSS.n1359 VSUBS 0.0148f
C1863 VSS.n1360 VSUBS 0.0129f
C1864 VSS.n1361 VSUBS 0.0189f
C1865 VSS.n1362 VSUBS 0.00845f
C1866 VSS.n1363 VSUBS 0.0149f
C1867 VSS.n1364 VSUBS 0.00483f
C1868 VSS.n1365 VSUBS 0.00411f
C1869 VSS.n1366 VSUBS 0.00895f
C1870 VSS.n1367 VSUBS 0.00774f
C1871 VSS.n1368 VSUBS 0.00629f
C1872 VSS.n1369 VSUBS 0.0148f
C1873 VSS.n1370 VSUBS 0.0253f
C1874 VSS.n1371 VSUBS 0.00646f
C1875 VSS.n1372 VSUBS 0.0169f
C1876 VSS.n1373 VSUBS 0.00677f
C1877 VSS.n1374 VSUBS 0.00314f
C1878 VSS.n1375 VSUBS 0.00339f
C1879 VSS.n1376 VSUBS 0.00596f
C1880 VSS.n1378 VSUBS 0.0163f
C1881 VSS.n1379 VSUBS 0.00497f
C1882 VSS.n1381 VSUBS 0.0148f
C1883 VSS.n1382 VSUBS 0.0224f
C1884 VSS.n1383 VSUBS 0.0109f
C1885 VSS.n1384 VSUBS 0.00774f
C1886 VSS.n1385 VSUBS 0.00339f
C1887 VSS.n1386 VSUBS 0.00314f
C1888 VSS.n1387 VSUBS 0.00646f
C1889 VSS.n1388 VSUBS 0.0169f
C1890 VSS.n1389 VSUBS 0.00774f
C1891 VSS.n1390 VSUBS 0.0109f
C1892 VSS.n1391 VSUBS 0.013f
C1893 VSS.n1392 VSUBS 0.0133f
C1894 VSS.n1393 VSUBS 0.0118f
C1895 VSS.n1394 VSUBS 0.00751f
C1896 VSS.n1395 VSUBS 0.0144f
C1897 VSS.n1396 VSUBS 0.0162f
C1898 VSS.n1397 VSUBS 0.00751f
C1899 VSS.n1398 VSUBS 0.0156f
C1900 VSS.n1399 VSUBS 0.015f
C1901 VSS.n1400 VSUBS 0.00751f
C1902 VSS.n1401 VSUBS 0.0118f
C1903 VSS.n1402 VSUBS 0.0127f
C1904 VSS.n1403 VSUBS 0.00664f
C1905 VSS.n1404 VSUBS 0.00693f
C1906 VSS.n1405 VSUBS 0.013f
C1907 VSS.n1406 VSUBS 0.0127f
C1908 VSS.n1407 VSUBS 0.00664f
C1909 VSS.n1408 VSUBS 0.00693f
C1910 VSS.n1409 VSUBS 0.013f
C1911 VSS.n1410 VSUBS 0.0116f
C1912 VSS.n1411 VSUBS 0.00751f
C1913 VSS.n1412 VSUBS 0.0153f
C1914 VSS.n1413 VSUBS 0.0153f
C1915 VSS.n1414 VSUBS 0.00751f
C1916 VSS.n1415 VSUBS 0.0165f
C1917 VSS.n1416 VSUBS 0.0142f
C1918 VSS.n1417 VSUBS 0.00751f
C1919 VSS.n1418 VSUBS 0.0121f
C1920 VSS.n1419 VSUBS 0.013f
C1921 VSS.t8 VSUBS 0.0256f
C1922 VSS.n1420 VSUBS 0.00596f
C1923 VSS.n1421 VSUBS 0.0148f
C1924 VSS.n1422 VSUBS 0.00497f
C1925 VSS.n1423 VSUBS 0.0148f
C1926 VSS.n1424 VSUBS 0.0253f
C1927 VSS.n1425 VSUBS 0.0109f
C1928 VSS.n1426 VSUBS 0.00677f
C1929 VSS.n1427 VSUBS 0.00629f
C1930 VSS.n1428 VSUBS 0.00798f
C1931 VSS.n1429 VSUBS 0.00871f
C1932 VSS.n1430 VSUBS 0.00411f
C1933 VSS.n1431 VSUBS 0.0209f
C1934 VSS.n1432 VSUBS 0.00745f
C1935 VSS.n1433 VSUBS 0.0148f
C1936 VSS.n1434 VSUBS 0.00298f
C1937 VSS.n1436 VSUBS 0.0148f
C1938 VSS.n1437 VSUBS 0.0253f
C1939 VSS.n1438 VSUBS 0.0109f
C1940 VSS.n1439 VSUBS 0.00484f
C1941 VSS.n1440 VSUBS 0.00629f
C1942 VSS.n1441 VSUBS 0.00895f
C1943 VSS.n1442 VSUBS 0.00967f
C1944 VSS.n1443 VSUBS 0.00411f
C1945 VSS.n1444 VSUBS 0.0229f
C1946 VSS.n1446 VSUBS 0.0402f
C1947 VSS.n1447 VSUBS 0.0163f
C1948 VSS.n1448 VSUBS 0.00845f
C1949 VSS.n1449 VSUBS 0.0109f
C1950 VSS.n1450 VSUBS 0.0029f
C1951 VSS.n1451 VSUBS 0.00459f
C1952 VSS.n1452 VSUBS 0.231f
C1953 VSS.n1453 VSUBS 0.00774f
C1954 VSS.n1454 VSUBS 0.0106f
C1955 VSS.n1455 VSUBS 0.0148f
C1956 VSS.n1456 VSUBS 0.0348f
C1957 VSS.n1458 VSUBS 0.0148f
C1958 VSS.n1459 VSUBS 0.0214f
C1959 VSS.n1460 VSUBS 0.0338f
C1960 VSS.n1461 VSUBS 0.00556f
C1961 VSS.n1462 VSUBS 0.00581f
C1962 VSS.n1463 VSUBS 0.0109f
C1963 VSS.n1464 VSUBS 0.0106f
C1964 VSS.n1465 VSUBS 0.00556f
C1965 VSS.n1466 VSUBS 0.0236f
C1966 VSS.n1467 VSUBS 0.0137f
C1967 VSS.n1468 VSUBS 0.0168f
C1968 VSS.n1469 VSUBS 0.0107f
C1969 VSS.n1470 VSUBS 0.0168f
C1970 VSS.n1471 VSUBS 0.0107f
C1971 VSS.n1472 VSUBS 0.0168f
C1972 VSS.n1473 VSUBS 0.0107f
C1973 VSS.n1474 VSUBS 0.0168f
C1974 VSS.n1475 VSUBS 0.0107f
C1975 VSS.n1476 VSUBS 0.0236f
C1976 VSS.n1477 VSUBS 0.0137f
C1977 VSS.n1478 VSUBS 0.0352f
C1978 VSS.n1480 VSUBS 0.0148f
C1979 VSS.n1481 VSUBS 0.0353f
C1980 VSS.n1482 VSUBS 0.0214f
C1981 VSS.n1483 VSUBS 0.00581f
C1982 VSS.n1484 VSUBS 0.0109f
C1983 VSS.n1485 VSUBS 0.00967f
C1984 VSS.n1486 VSUBS 0.00629f
C1985 VSS.n1487 VSUBS 0.0263f
C1986 VSS.n1488 VSUBS 0.0163f
C1987 VSS.n1489 VSUBS 0.00298f
C1988 VSS.n1490 VSUBS 0.0148f
C1989 VSS.n1491 VSUBS 0.00696f
C1990 VSS.n1492 VSUBS 0.00546f
C1991 VSS.n1493 VSUBS 0.0288f
C1992 VSS.n1494 VSUBS 0.0029f
C1993 VSS.n1495 VSUBS 0.00411f
C1994 VSS.n1496 VSUBS 0.00992f
C1995 VSS.n1497 VSUBS 0.00871f
C1996 VSS.n1498 VSUBS 0.00629f
C1997 VSS.n1499 VSUBS 0.0263f
C1998 VSS.n1501 VSUBS 0.0148f
C1999 VSS.n1502 VSUBS 0.00298f
C2000 VSS.n1503 VSUBS 0.0148f
C2001 VSS.n1504 VSUBS 0.00497f
C2002 VSS.n1505 VSUBS 0.00546f
C2003 VSS.n1506 VSUBS 0.0278f
C2004 VSS.n1507 VSUBS 0.00483f
C2005 VSS.n1508 VSUBS 0.00411f
C2006 VSS.n1509 VSUBS 0.00895f
C2007 VSS.n1510 VSUBS 0.00774f
C2008 VSS.n1511 VSUBS 0.00629f
C2009 VSS.n1513 VSUBS 0.0148f
C2010 VSS.n1514 VSUBS 0.00199f
C2011 VSS.n1515 VSUBS 0.00546f
C2012 VSS.n1516 VSUBS 0.0298f
C2013 VSS.n1517 VSUBS 0.00677f
C2014 VSS.n1518 VSUBS 0.00314f
C2015 VSS.n1519 VSUBS 0.00339f
C2016 VSS.n1520 VSUBS 0.00199f
C2017 VSS.n1522 VSUBS 0.0148f
C2018 VSS.n1523 VSUBS 0.00497f
C2019 VSS.n1524 VSUBS 0.0263f
C2020 VSS.n1525 VSUBS 0.00774f
C2021 VSS.n1526 VSUBS 0.00339f
C2022 VSS.n1527 VSUBS 0.00314f
C2023 VSS.n1529 VSUBS 0.0148f
C2024 VSS.n1530 VSUBS 0.00199f
C2025 VSS.n1531 VSUBS 0.00546f
C2026 VSS.n1532 VSUBS 0.0268f
C2027 VSS.n1533 VSUBS 0.00774f
C2028 VSS.n1534 VSUBS 0.0109f
C2029 VSS.n1535 VSUBS 0.013f
C2030 VSS.n1536 VSUBS 0.0133f
C2031 VSS.n1537 VSUBS 0.0118f
C2032 VSS.n1538 VSUBS 0.00751f
C2033 VSS.n1539 VSUBS 0.0144f
C2034 VSS.n1540 VSUBS 0.0162f
C2035 VSS.n1541 VSUBS 0.00751f
C2036 VSS.n1542 VSUBS 0.0156f
C2037 VSS.n1543 VSUBS 0.015f
C2038 VSS.n1544 VSUBS 0.00751f
C2039 VSS.n1545 VSUBS 0.0118f
C2040 VSS.n1546 VSUBS 0.0127f
C2041 VSS.n1547 VSUBS 0.00664f
C2042 VSS.n1548 VSUBS 0.00693f
C2043 VSS.n1549 VSUBS 0.013f
C2044 VSS.n1550 VSUBS 0.0127f
C2045 VSS.n1551 VSUBS 0.00664f
C2046 VSS.n1552 VSUBS 0.00693f
C2047 VSS.n1553 VSUBS 0.013f
C2048 VSS.n1554 VSUBS 0.0116f
C2049 VSS.n1555 VSUBS 0.00751f
C2050 VSS.n1556 VSUBS 0.0153f
C2051 VSS.n1557 VSUBS 0.0153f
C2052 VSS.n1558 VSUBS 0.00751f
C2053 VSS.n1559 VSUBS 0.0165f
C2054 VSS.n1560 VSUBS 0.0142f
C2055 VSS.n1561 VSUBS 0.00751f
C2056 VSS.n1562 VSUBS 0.0121f
C2057 VSS.n1563 VSUBS 0.013f
C2058 VSS.n1564 VSUBS 0.00199f
C2059 VSS.n1565 VSUBS 0.0163f
C2060 VSS.n1566 VSUBS 0.00497f
C2061 VSS.n1567 VSUBS 0.0293f
C2062 VSS.n1568 VSUBS 0.00677f
C2063 VSS.n1569 VSUBS 0.00629f
C2064 VSS.n1570 VSUBS 0.00798f
C2065 VSS.n1571 VSUBS 0.00871f
C2066 VSS.n1572 VSUBS 0.00411f
C2067 VSS.n1573 VSUBS 0.0278f
C2068 VSS.n1574 VSUBS 0.0148f
C2069 VSS.n1575 VSUBS 0.00546f
C2070 VSS.n1576 VSUBS 0.00596f
C2071 VSS.n1577 VSUBS 0.0224f
C2072 VSS.n1578 VSUBS 0.00484f
C2073 VSS.n1579 VSUBS 0.00629f
C2074 VSS.n1580 VSUBS 0.00895f
C2075 VSS.n1581 VSUBS 0.00967f
C2076 VSS.n1582 VSUBS 0.00411f
C2077 VSS.n1583 VSUBS 0.0168f
C2078 VSS.n1584 VSUBS 0.0107f
C2079 VSS.n1585 VSUBS 0.0168f
C2080 VSS.n1586 VSUBS 0.0107f
C2081 VSS.n1587 VSUBS 0.0168f
C2082 VSS.n1588 VSUBS 0.0107f
C2083 VSS.n1589 VSUBS 0.0168f
C2084 VSS.n1590 VSUBS 0.0107f
C2085 VSS.n1591 VSUBS 0.0236f
C2086 VSS.n1592 VSUBS 0.0137f
C2087 VSS.n1593 VSUBS 0.0337f
C2088 VSS.n1594 VSUBS 0.00845f
C2089 VSS.n1595 VSUBS 0.0148f
C2090 VSS.n1596 VSUBS 0.00745f
C2091 VSS.n1597 VSUBS 0.00596f
C2092 VSS.n1598 VSUBS 0.0288f
C2093 VSS.n1599 VSUBS 0.0029f
C2094 VSS.n1600 VSUBS 0.00629f
C2095 VSS.n1601 VSUBS 0.00992f
C2096 VSS.n1602 VSUBS 0.0106f
C2097 VSS.n1604 VSUBS 0.0148f
C2098 VSS.n1605 VSUBS 0.0348f
C2099 VSS.n1606 VSUBS 0.0402f
C2100 VSS.n1607 VSUBS 0.0163f
C2101 VSS.n1608 VSUBS 0.0268f
C2102 VSS.n1609 VSUBS 0.0149f
C2103 VSS.n1610 VSUBS 0.00556f
C2104 VSS.n1611 VSUBS 0.00581f
C2105 VSS.n1612 VSUBS 0.0109f
C2106 VSS.n1613 VSUBS 0.0106f
C2107 VSS.n1614 VSUBS 0.00556f
C2108 VSS.n1616 VSUBS 0.0148f
C2109 VSS.n1617 VSUBS 0.0278f
C2110 VSS.n1618 VSUBS 0.0148f
C2111 VSS.n1619 VSUBS 0.0293f
C2112 VSS.n1620 VSUBS 2.92f
C2113 VSS.n1621 VSUBS 1.55f
C2114 VSS.n1623 VSUBS 0.0148f
C2115 VSS.n1624 VSUBS 0.0248f
C2116 VSS.n1625 VSUBS 0.0149f
C2117 VSS.n1626 VSUBS 0.00581f
C2118 VSS.n1627 VSUBS 0.0109f
C2119 VSS.n1628 VSUBS 0.00967f
C2120 VSS.n1629 VSUBS 0.00629f
C2121 VSS.n1630 VSUBS 0.0189f
C2122 VSS.n1631 VSUBS 0.0148f
C2123 VSS.n1632 VSUBS 0.00795f
C2124 VSS.n1633 VSUBS 0.00447f
C2125 VSS.n1634 VSUBS 0.0109f
C2126 VSS.n1635 VSUBS 0.0029f
C2127 VSS.n1636 VSUBS 0.00411f
C2128 VSS.n1637 VSUBS 0.00992f
C2129 VSS.n1638 VSUBS 0.00871f
C2130 VSS.n1639 VSUBS 0.00629f
C2131 VSS.n1640 VSUBS 0.0148f
C2132 VSS.n1641 VSUBS 0.0253f
C2133 VSS.n1642 VSUBS 0.0189f
C2134 VSS.n1644 VSUBS 0.0326f
C2135 VSS.n1645 VSUBS 0.00596f
C2136 VSS.n1646 VSUBS 0.00447f
C2137 VSS.n1647 VSUBS 0.0129f
C2138 VSS.n1648 VSUBS 0.00483f
C2139 VSS.n1649 VSUBS 0.00411f
C2140 VSS.n1650 VSUBS 0.00895f
C2141 VSS.n1651 VSUBS 0.00774f
C2142 VSS.n1652 VSUBS 0.00629f
C2143 VSS.n1654 VSUBS 0.0148f
C2144 VSS.n1655 VSUBS 0.0253f
C2145 VSS.n1656 VSUBS 0.00646f
C2146 VSS.n1657 VSUBS 0.0149f
C2147 VSS.n1658 VSUBS 0.00677f
C2148 VSS.n1659 VSUBS 0.00314f
C2149 VSS.n1660 VSUBS 0.00339f
C2150 VSS.n1661 VSUBS 0.00696f
C2151 VSS.n1662 VSUBS 0.0169f
C2152 VSS.n1663 VSUBS 0.00774f
C2153 VSS.n1664 VSUBS 0.00992f
C2154 VSS.n1665 VSUBS 0.00629f
C2155 VSS.n1666 VSUBS 0.0029f
C2156 VSS.n1667 VSUBS 0.00411f
C2157 VSS.n1668 VSUBS 0.00967f
C2158 VSS.n1669 VSUBS 0.00895f
C2159 VSS.n1670 VSUBS 0.00629f
C2160 VSS.n1671 VSUBS 0.00484f
C2161 VSS.n1672 VSUBS 0.00411f
C2162 VSS.n1673 VSUBS 0.00871f
C2163 VSS.n1674 VSUBS 0.00798f
C2164 VSS.n1675 VSUBS 0.00629f
C2165 VSS.n1676 VSUBS 0.00677f
C2166 VSS.n1677 VSUBS 0.00339f
C2167 VSS.n1678 VSUBS 0.00314f
C2168 VSS.n1679 VSUBS 0.00774f
C2169 VSS.n1680 VSUBS 0.0109f
C2170 VSS.n1681 VSUBS 0.013f
C2171 VSS.n1682 VSUBS 0.0133f
C2172 VSS.n1683 VSUBS 0.0118f
C2173 VSS.n1684 VSUBS 0.00751f
C2174 VSS.n1685 VSUBS 0.0144f
C2175 VSS.n1686 VSUBS 0.0162f
C2176 VSS.n1687 VSUBS 0.00751f
C2177 VSS.n1688 VSUBS 0.0156f
C2178 VSS.n1689 VSUBS 0.015f
C2179 VSS.n1690 VSUBS 0.00751f
C2180 VSS.n1691 VSUBS 0.0118f
C2181 VSS.n1692 VSUBS 0.0127f
C2182 VSS.n1693 VSUBS 0.00664f
C2183 VSS.n1694 VSUBS 0.0106f
C2184 VSS.n1695 VSUBS 0.00556f
C2185 VSS.n1696 VSUBS 0.00581f
C2186 VSS.n1697 VSUBS 0.00693f
C2187 VSS.n1698 VSUBS 0.013f
C2188 VSS.n1699 VSUBS 0.0127f
C2189 VSS.n1700 VSUBS 0.0109f
C2190 VSS.n1701 VSUBS 0.0106f
C2191 VSS.n1702 VSUBS 0.0357f
C2192 VSS.n1703 VSUBS 0.00556f
C2193 VSS.n1704 VSUBS 0.0117f
C2194 VSS.n1705 VSUBS 0.139f
C2195 VSS.n1706 VSUBS 0.0204f
C2196 VSS.t39 VSUBS 0.0109f
C2197 VSS.t48 VSUBS 0.0109f
C2198 VSS.n1707 VSUBS 0.0263f
C2199 VSS.n1708 VSUBS 0.00951f
C2200 VSS.n1709 VSUBS 0.0254f
C2201 VSS.n1710 VSUBS 0.00679f
C2202 VSS.n1711 VSUBS 0.00335f
C2203 VSS.n1712 VSUBS 0.0107f
C2204 VSS.n1713 VSUBS 0.199f
C2205 VSS.n1714 VSUBS 0.0837f
C2206 VSS.n1715 VSUBS 0.0174f
C2207 VSS.t112 VSUBS 0.0109f
C2208 VSS.t29 VSUBS 0.0109f
C2209 VSS.n1716 VSUBS 0.0263f
C2210 VSS.n1717 VSUBS 0.00951f
C2211 VSS.n1718 VSUBS 0.0254f
C2212 VSS.n1719 VSUBS 0.00679f
C2213 VSS.n1720 VSUBS 0.00335f
C2214 VSS.n1721 VSUBS 0.0107f
C2215 VSS.n1722 VSUBS 0.0816f
C2216 VSS.n1723 VSUBS 0.0837f
C2217 VSS.n1724 VSUBS 0.0174f
C2218 VSS.t42 VSUBS 0.0109f
C2219 VSS.t84 VSUBS 0.0109f
C2220 VSS.n1725 VSUBS 0.0263f
C2221 VSS.n1726 VSUBS 0.00951f
C2222 VSS.n1727 VSUBS 0.0254f
C2223 VSS.n1728 VSUBS 0.00679f
C2224 VSS.n1729 VSUBS 0.00335f
C2225 VSS.n1730 VSUBS 0.0107f
C2226 VSS.n1731 VSUBS 0.0816f
C2227 VSS.n1732 VSUBS 0.0837f
C2228 VSS.n1733 VSUBS 0.0174f
C2229 VSS.t89 VSUBS 0.0109f
C2230 VSS.t55 VSUBS 0.0109f
C2231 VSS.n1734 VSUBS 0.0263f
C2232 VSS.n1735 VSUBS 0.00951f
C2233 VSS.n1736 VSUBS 0.0254f
C2234 VSS.n1737 VSUBS 0.00679f
C2235 VSS.n1738 VSUBS 0.00335f
C2236 VSS.n1739 VSUBS 0.0107f
C2237 VSS.n1740 VSUBS 0.0816f
C2238 VSS.n1741 VSUBS 0.0837f
C2239 VSS.n1742 VSUBS 0.0174f
C2240 VSS.t27 VSUBS 0.0109f
C2241 VSS.t78 VSUBS 0.0109f
C2242 VSS.n1743 VSUBS 0.0263f
C2243 VSS.n1744 VSUBS 0.00951f
C2244 VSS.n1745 VSUBS 0.0254f
C2245 VSS.n1746 VSUBS 0.00679f
C2246 VSS.n1747 VSUBS 0.00335f
C2247 VSS.n1748 VSUBS 0.0107f
C2248 VSS.n1749 VSUBS 0.0816f
C2249 VSS.n1750 VSUBS 0.0837f
C2250 VSS.n1751 VSUBS 0.0174f
C2251 VSS.t131 VSUBS 0.0109f
C2252 VSS.t136 VSUBS 0.0109f
C2253 VSS.n1752 VSUBS 0.0263f
C2254 VSS.n1753 VSUBS 0.00951f
C2255 VSS.n1754 VSUBS 0.0254f
C2256 VSS.n1755 VSUBS 0.00679f
C2257 VSS.n1756 VSUBS 0.00335f
C2258 VSS.n1757 VSUBS 0.0107f
C2259 VSS.n1758 VSUBS 0.0816f
C2260 VSS.n1759 VSUBS 0.0837f
C2261 VSS.n1760 VSUBS 0.0174f
C2262 VSS.t86 VSUBS 0.0109f
C2263 VSS.t93 VSUBS 0.0109f
C2264 VSS.n1761 VSUBS 0.0263f
C2265 VSS.n1762 VSUBS 0.00951f
C2266 VSS.n1763 VSUBS 0.0254f
C2267 VSS.n1764 VSUBS 0.00679f
C2268 VSS.n1765 VSUBS 0.00335f
C2269 VSS.n1766 VSUBS 0.0107f
C2270 VSS.n1767 VSUBS 0.0816f
C2271 VSS.n1768 VSUBS 0.0837f
C2272 VSS.n1769 VSUBS 0.0174f
C2273 VSS.t132 VSUBS 0.0109f
C2274 VSS.t123 VSUBS 0.0109f
C2275 VSS.n1770 VSUBS 0.0263f
C2276 VSS.n1771 VSUBS 0.00951f
C2277 VSS.n1772 VSUBS 0.0254f
C2278 VSS.n1773 VSUBS 0.00679f
C2279 VSS.n1774 VSUBS 0.00335f
C2280 VSS.n1775 VSUBS 0.0107f
C2281 VSS.n1776 VSUBS 0.0816f
C2282 VSS.n1777 VSUBS 0.0837f
C2283 VSS.n1778 VSUBS 0.0174f
C2284 VSS.t110 VSUBS 0.0109f
C2285 VSS.t25 VSUBS 0.0109f
C2286 VSS.n1779 VSUBS 0.0263f
C2287 VSS.n1780 VSUBS 0.00951f
C2288 VSS.n1781 VSUBS 0.0254f
C2289 VSS.n1782 VSUBS 0.00679f
C2290 VSS.n1783 VSUBS 0.00335f
C2291 VSS.n1784 VSUBS 0.0107f
C2292 VSS.n1785 VSUBS 0.0816f
C2293 VSS.n1786 VSUBS 0.0837f
C2294 VSS.n1787 VSUBS 0.0174f
C2295 VSS.t19 VSUBS 0.0109f
C2296 VSS.t98 VSUBS 0.0109f
C2297 VSS.n1788 VSUBS 0.0263f
C2298 VSS.n1789 VSUBS 0.00951f
C2299 VSS.n1790 VSUBS 0.0254f
C2300 VSS.n1791 VSUBS 0.00679f
C2301 VSS.n1792 VSUBS 0.00335f
C2302 VSS.n1793 VSUBS 0.0107f
C2303 VSS.n1794 VSUBS 0.0816f
C2304 VSS.n1795 VSUBS 0.0837f
C2305 VSS.n1796 VSUBS 0.0174f
C2306 VSS.t88 VSUBS 0.0109f
C2307 VSS.t53 VSUBS 0.0109f
C2308 VSS.n1797 VSUBS 0.0263f
C2309 VSS.n1798 VSUBS 0.00951f
C2310 VSS.n1799 VSUBS 0.0254f
C2311 VSS.n1800 VSUBS 0.00679f
C2312 VSS.n1801 VSUBS 0.00335f
C2313 VSS.n1802 VSUBS 0.0107f
C2314 VSS.n1803 VSUBS 0.0816f
C2315 VSS.n1804 VSUBS 0.0837f
C2316 VSS.n1805 VSUBS 0.0174f
C2317 VSS.t87 VSUBS 0.0109f
C2318 VSS.t83 VSUBS 0.0109f
C2319 VSS.n1806 VSUBS 0.0263f
C2320 VSS.n1807 VSUBS 0.00951f
C2321 VSS.n1808 VSUBS 0.0254f
C2322 VSS.n1809 VSUBS 0.00679f
C2323 VSS.n1810 VSUBS 0.00335f
C2324 VSS.n1811 VSUBS 0.0107f
C2325 VSS.n1812 VSUBS 0.0816f
C2326 VSS.n1813 VSUBS 0.0837f
C2327 VSS.n1814 VSUBS 0.0174f
C2328 VSS.t40 VSUBS 0.0109f
C2329 VSS.t28 VSUBS 0.0109f
C2330 VSS.n1815 VSUBS 0.0263f
C2331 VSS.n1816 VSUBS 0.00951f
C2332 VSS.n1817 VSUBS 0.0254f
C2333 VSS.n1818 VSUBS 0.00679f
C2334 VSS.n1819 VSUBS 0.00335f
C2335 VSS.n1820 VSUBS 0.0107f
C2336 VSS.n1821 VSUBS 0.0816f
C2337 VSS.n1822 VSUBS 0.0837f
C2338 VSS.n1823 VSUBS 0.0174f
C2339 VSS.t109 VSUBS 0.0109f
C2340 VSS.t81 VSUBS 0.0109f
C2341 VSS.n1824 VSUBS 0.0263f
C2342 VSS.n1825 VSUBS 0.00951f
C2343 VSS.n1826 VSUBS 0.0254f
C2344 VSS.n1827 VSUBS 0.00679f
C2345 VSS.n1828 VSUBS 0.00335f
C2346 VSS.n1829 VSUBS 0.0107f
C2347 VSS.n1830 VSUBS 0.0816f
C2348 VSS.n1831 VSUBS 0.0837f
C2349 VSS.n1832 VSUBS 0.0174f
C2350 VSS.t36 VSUBS 0.0109f
C2351 VSS.t118 VSUBS 0.0109f
C2352 VSS.n1833 VSUBS 0.0263f
C2353 VSS.n1834 VSUBS 0.00951f
C2354 VSS.n1835 VSUBS 0.0254f
C2355 VSS.n1836 VSUBS 0.00679f
C2356 VSS.n1837 VSUBS 0.00335f
C2357 VSS.n1838 VSUBS 0.0107f
C2358 VSS.n1839 VSUBS 0.0816f
C2359 VSS.n1840 VSUBS 0.0837f
C2360 VSS.n1841 VSUBS 0.0174f
C2361 VSS.t107 VSUBS 0.0109f
C2362 VSS.t65 VSUBS 0.0109f
C2363 VSS.n1842 VSUBS 0.0263f
C2364 VSS.n1843 VSUBS 0.00951f
C2365 VSS.n1844 VSUBS 0.0254f
C2366 VSS.n1845 VSUBS 0.00679f
C2367 VSS.n1846 VSUBS 0.00335f
C2368 VSS.n1847 VSUBS 0.0107f
C2369 VSS.n1848 VSUBS 0.0816f
C2370 VSS.n1849 VSUBS 0.0837f
C2371 VSS.n1850 VSUBS 0.0174f
C2372 VSS.t16 VSUBS 0.0109f
C2373 VSS.t114 VSUBS 0.0109f
C2374 VSS.n1851 VSUBS 0.0263f
C2375 VSS.n1852 VSUBS 0.00951f
C2376 VSS.n1853 VSUBS 0.0254f
C2377 VSS.n1854 VSUBS 0.00679f
C2378 VSS.n1855 VSUBS 0.00335f
C2379 VSS.n1856 VSUBS 0.0107f
C2380 VSS.n1857 VSUBS 0.0816f
C2381 VSS.n1858 VSUBS 0.0837f
C2382 VSS.n1859 VSUBS 0.0174f
C2383 VSS.t70 VSUBS 0.0109f
C2384 VSS.t62 VSUBS 0.0109f
C2385 VSS.n1860 VSUBS 0.0263f
C2386 VSS.n1861 VSUBS 0.00951f
C2387 VSS.n1862 VSUBS 0.0254f
C2388 VSS.n1863 VSUBS 0.00679f
C2389 VSS.n1864 VSUBS 0.00335f
C2390 VSS.n1865 VSUBS 0.0107f
C2391 VSS.n1866 VSUBS 0.0816f
C2392 VSS.n1867 VSUBS 0.0837f
C2393 VSS.n1868 VSUBS 0.0174f
C2394 VSS.t135 VSUBS 0.0109f
C2395 VSS.t91 VSUBS 0.0109f
C2396 VSS.n1869 VSUBS 0.0263f
C2397 VSS.n1870 VSUBS 0.00951f
C2398 VSS.n1871 VSUBS 0.0254f
C2399 VSS.n1872 VSUBS 0.00679f
C2400 VSS.n1873 VSUBS 0.00335f
C2401 VSS.n1874 VSUBS 0.0107f
C2402 VSS.n1875 VSUBS 0.0816f
C2403 VSS.n1876 VSUBS 0.0837f
C2404 VSS.n1877 VSUBS 0.0174f
C2405 VSS.t51 VSUBS 0.0109f
C2406 VSS.t43 VSUBS 0.0109f
C2407 VSS.n1878 VSUBS 0.0263f
C2408 VSS.n1879 VSUBS 0.00951f
C2409 VSS.n1880 VSUBS 0.0254f
C2410 VSS.n1881 VSUBS 0.00679f
C2411 VSS.n1882 VSUBS 0.00335f
C2412 VSS.n1883 VSUBS 0.0107f
C2413 VSS.n1884 VSUBS 0.0782f
C2414 VSS.n1885 VSUBS 0.0204f
C2415 VSS.t101 VSUBS 0.0109f
C2416 VSS.t111 VSUBS 0.0109f
C2417 VSS.n1886 VSUBS 0.0263f
C2418 VSS.n1887 VSUBS 0.00951f
C2419 VSS.n1888 VSUBS 0.0254f
C2420 VSS.n1889 VSUBS 0.00679f
C2421 VSS.n1890 VSUBS 0.00335f
C2422 VSS.n1891 VSUBS 0.0107f
C2423 VSS.n1892 VSUBS 0.199f
C2424 VSS.n1893 VSUBS 0.0837f
C2425 VSS.n1894 VSUBS 0.0174f
C2426 VSS.t58 VSUBS 0.0109f
C2427 VSS.t97 VSUBS 0.0109f
C2428 VSS.n1895 VSUBS 0.0263f
C2429 VSS.n1896 VSUBS 0.00951f
C2430 VSS.n1897 VSUBS 0.0254f
C2431 VSS.n1898 VSUBS 0.00679f
C2432 VSS.n1899 VSUBS 0.00335f
C2433 VSS.n1900 VSUBS 0.0107f
C2434 VSS.n1901 VSUBS 0.0816f
C2435 VSS.n1902 VSUBS 0.0837f
C2436 VSS.n1903 VSUBS 0.0174f
C2437 VSS.t103 VSUBS 0.0109f
C2438 VSS.t22 VSUBS 0.0109f
C2439 VSS.n1904 VSUBS 0.0263f
C2440 VSS.n1905 VSUBS 0.00951f
C2441 VSS.n1906 VSUBS 0.0254f
C2442 VSS.n1907 VSUBS 0.00679f
C2443 VSS.n1908 VSUBS 0.00335f
C2444 VSS.n1909 VSUBS 0.0107f
C2445 VSS.n1910 VSUBS 0.0816f
C2446 VSS.n1911 VSUBS 0.0837f
C2447 VSS.n1912 VSUBS 0.0174f
C2448 VSS.t33 VSUBS 0.0109f
C2449 VSS.t122 VSUBS 0.0109f
C2450 VSS.n1913 VSUBS 0.0263f
C2451 VSS.n1914 VSUBS 0.00951f
C2452 VSS.n1915 VSUBS 0.0254f
C2453 VSS.n1916 VSUBS 0.00679f
C2454 VSS.n1917 VSUBS 0.00335f
C2455 VSS.n1918 VSUBS 0.0107f
C2456 VSS.n1919 VSUBS 0.0816f
C2457 VSS.n1920 VSUBS 0.0837f
C2458 VSS.n1921 VSUBS 0.0174f
C2459 VSS.t95 VSUBS 0.0109f
C2460 VSS.t18 VSUBS 0.0109f
C2461 VSS.n1922 VSUBS 0.0263f
C2462 VSS.n1923 VSUBS 0.00951f
C2463 VSS.n1924 VSUBS 0.0254f
C2464 VSS.n1925 VSUBS 0.00679f
C2465 VSS.n1926 VSUBS 0.00335f
C2466 VSS.n1927 VSUBS 0.0107f
C2467 VSS.n1928 VSUBS 0.0816f
C2468 VSS.n1929 VSUBS 0.0837f
C2469 VSS.n1930 VSUBS 0.0174f
C2470 VSS.t72 VSUBS 0.0109f
C2471 VSS.t75 VSUBS 0.0109f
C2472 VSS.n1931 VSUBS 0.0263f
C2473 VSS.n1932 VSUBS 0.00951f
C2474 VSS.n1933 VSUBS 0.0254f
C2475 VSS.n1934 VSUBS 0.00679f
C2476 VSS.n1935 VSUBS 0.00335f
C2477 VSS.n1936 VSUBS 0.0107f
C2478 VSS.n1937 VSUBS 0.0816f
C2479 VSS.n1938 VSUBS 0.0837f
C2480 VSS.n1939 VSUBS 0.0174f
C2481 VSS.t26 VSUBS 0.0109f
C2482 VSS.t38 VSUBS 0.0109f
C2483 VSS.n1940 VSUBS 0.0263f
C2484 VSS.n1941 VSUBS 0.00951f
C2485 VSS.n1942 VSUBS 0.0254f
C2486 VSS.n1943 VSUBS 0.00679f
C2487 VSS.n1944 VSUBS 0.00335f
C2488 VSS.n1945 VSUBS 0.0107f
C2489 VSS.n1946 VSUBS 0.0816f
C2490 VSS.n1947 VSUBS 0.0837f
C2491 VSS.n1948 VSUBS 0.0174f
C2492 VSS.t73 VSUBS 0.0109f
C2493 VSS.t63 VSUBS 0.0109f
C2494 VSS.n1949 VSUBS 0.0263f
C2495 VSS.n1950 VSUBS 0.00951f
C2496 VSS.n1951 VSUBS 0.0254f
C2497 VSS.n1952 VSUBS 0.00679f
C2498 VSS.n1953 VSUBS 0.00335f
C2499 VSS.n1954 VSUBS 0.0107f
C2500 VSS.n1955 VSUBS 0.0816f
C2501 VSS.n1956 VSUBS 0.0837f
C2502 VSS.n1957 VSUBS 0.0174f
C2503 VSS.t57 VSUBS 0.0109f
C2504 VSS.t92 VSUBS 0.0109f
C2505 VSS.n1958 VSUBS 0.0263f
C2506 VSS.n1959 VSUBS 0.00951f
C2507 VSS.n1960 VSUBS 0.0254f
C2508 VSS.n1961 VSUBS 0.00679f
C2509 VSS.n1962 VSUBS 0.00335f
C2510 VSS.n1963 VSUBS 0.0107f
C2511 VSS.n1964 VSUBS 0.0816f
C2512 VSS.n1965 VSUBS 0.0837f
C2513 VSS.n1966 VSUBS 0.0174f
C2514 VSS.t85 VSUBS 0.0109f
C2515 VSS.t44 VSUBS 0.0109f
C2516 VSS.n1967 VSUBS 0.0263f
C2517 VSS.n1968 VSUBS 0.00951f
C2518 VSS.n1969 VSUBS 0.0254f
C2519 VSS.n1970 VSUBS 0.00679f
C2520 VSS.n1971 VSUBS 0.00335f
C2521 VSS.n1972 VSUBS 0.0107f
C2522 VSS.n1973 VSUBS 0.0816f
C2523 VSS.n1974 VSUBS 0.0837f
C2524 VSS.n1975 VSUBS 0.0174f
C2525 VSS.t32 VSUBS 0.0109f
C2526 VSS.t120 VSUBS 0.0109f
C2527 VSS.n1976 VSUBS 0.0263f
C2528 VSS.n1977 VSUBS 0.00951f
C2529 VSS.n1978 VSUBS 0.0254f
C2530 VSS.n1979 VSUBS 0.00679f
C2531 VSS.n1980 VSUBS 0.00335f
C2532 VSS.n1981 VSUBS 0.0107f
C2533 VSS.n1982 VSUBS 0.0816f
C2534 VSS.n1983 VSUBS 0.0837f
C2535 VSS.n1984 VSUBS 0.0174f
C2536 VSS.t30 VSUBS 0.0109f
C2537 VSS.t21 VSUBS 0.0109f
C2538 VSS.n1985 VSUBS 0.0263f
C2539 VSS.n1986 VSUBS 0.00951f
C2540 VSS.n1987 VSUBS 0.0254f
C2541 VSS.n1988 VSUBS 0.00679f
C2542 VSS.n1989 VSUBS 0.00335f
C2543 VSS.n1990 VSUBS 0.0107f
C2544 VSS.n1991 VSUBS 0.0816f
C2545 VSS.n1992 VSUBS 0.0837f
C2546 VSS.n1993 VSUBS 0.0174f
C2547 VSS.t102 VSUBS 0.0109f
C2548 VSS.t96 VSUBS 0.0109f
C2549 VSS.n1994 VSUBS 0.0263f
C2550 VSS.n1995 VSUBS 0.00951f
C2551 VSS.n1996 VSUBS 0.0254f
C2552 VSS.n1997 VSUBS 0.00679f
C2553 VSS.n1998 VSUBS 0.00335f
C2554 VSS.n1999 VSUBS 0.0107f
C2555 VSS.n2000 VSUBS 0.0816f
C2556 VSS.n2001 VSUBS 0.0837f
C2557 VSS.n2002 VSUBS 0.0174f
C2558 VSS.t56 VSUBS 0.0109f
C2559 VSS.t20 VSUBS 0.0109f
C2560 VSS.n2003 VSUBS 0.0263f
C2561 VSS.n2004 VSUBS 0.00951f
C2562 VSS.n2005 VSUBS 0.0254f
C2563 VSS.n2006 VSUBS 0.00679f
C2564 VSS.n2007 VSUBS 0.00335f
C2565 VSS.n2008 VSUBS 0.0107f
C2566 VSS.n2009 VSUBS 0.0816f
C2567 VSS.n2010 VSUBS 0.0837f
C2568 VSS.n2011 VSUBS 0.0174f
C2569 VSS.t99 VSUBS 0.0109f
C2570 VSS.t60 VSUBS 0.0109f
C2571 VSS.n2012 VSUBS 0.0263f
C2572 VSS.n2013 VSUBS 0.00951f
C2573 VSS.n2014 VSUBS 0.0254f
C2574 VSS.n2015 VSUBS 0.00679f
C2575 VSS.n2016 VSUBS 0.00335f
C2576 VSS.n2017 VSUBS 0.0107f
C2577 VSS.n2018 VSUBS 0.0816f
C2578 VSS.n2019 VSUBS 0.0837f
C2579 VSS.n2020 VSUBS 0.0174f
C2580 VSS.t52 VSUBS 0.0109f
C2581 VSS.t129 VSUBS 0.0109f
C2582 VSS.n2021 VSUBS 0.0263f
C2583 VSS.n2022 VSUBS 0.00951f
C2584 VSS.n2023 VSUBS 0.0254f
C2585 VSS.n2024 VSUBS 0.00679f
C2586 VSS.n2025 VSUBS 0.00335f
C2587 VSS.n2026 VSUBS 0.0107f
C2588 VSS.n2027 VSUBS 0.0816f
C2589 VSS.n2028 VSUBS 0.0837f
C2590 VSS.n2029 VSUBS 0.0174f
C2591 VSS.t82 VSUBS 0.0109f
C2592 VSS.t59 VSUBS 0.0109f
C2593 VSS.n2030 VSUBS 0.0263f
C2594 VSS.n2031 VSUBS 0.00951f
C2595 VSS.n2032 VSUBS 0.0254f
C2596 VSS.n2033 VSUBS 0.00679f
C2597 VSS.n2034 VSUBS 0.00335f
C2598 VSS.n2035 VSUBS 0.0107f
C2599 VSS.n2036 VSUBS 0.0816f
C2600 VSS.n2037 VSUBS 0.0837f
C2601 VSS.n2038 VSUBS 0.0174f
C2602 VSS.t130 VSUBS 0.0109f
C2603 VSS.t127 VSUBS 0.0109f
C2604 VSS.n2039 VSUBS 0.0263f
C2605 VSS.n2040 VSUBS 0.00951f
C2606 VSS.n2041 VSUBS 0.0254f
C2607 VSS.n2042 VSUBS 0.00679f
C2608 VSS.n2043 VSUBS 0.00335f
C2609 VSS.n2044 VSUBS 0.0107f
C2610 VSS.n2045 VSUBS 0.0816f
C2611 VSS.n2046 VSUBS 0.0837f
C2612 VSS.n2047 VSUBS 0.0174f
C2613 VSS.t74 VSUBS 0.0109f
C2614 VSS.t35 VSUBS 0.0109f
C2615 VSS.n2048 VSUBS 0.0263f
C2616 VSS.n2049 VSUBS 0.00951f
C2617 VSS.n2050 VSUBS 0.0254f
C2618 VSS.n2051 VSUBS 0.00679f
C2619 VSS.n2052 VSUBS 0.00335f
C2620 VSS.n2053 VSUBS 0.0107f
C2621 VSS.n2054 VSUBS 0.0816f
C2622 VSS.n2055 VSUBS 0.0837f
C2623 VSS.n2056 VSUBS 0.0174f
C2624 VSS.t117 VSUBS 0.0109f
C2625 VSS.t106 VSUBS 0.0109f
C2626 VSS.n2057 VSUBS 0.0263f
C2627 VSS.n2058 VSUBS 0.00951f
C2628 VSS.n2059 VSUBS 0.0254f
C2629 VSS.n2060 VSUBS 0.00679f
C2630 VSS.n2061 VSUBS 0.00335f
C2631 VSS.n2062 VSUBS 0.0107f
C2632 VSS.n2063 VSUBS 0.0782f
C2633 VSS.n2064 VSUBS 0.0204f
C2634 VSS.t115 VSUBS 0.0109f
C2635 VSS.t124 VSUBS 0.0109f
C2636 VSS.n2065 VSUBS 0.0263f
C2637 VSS.n2066 VSUBS 0.00951f
C2638 VSS.n2067 VSUBS 0.0254f
C2639 VSS.n2068 VSUBS 0.00679f
C2640 VSS.n2069 VSUBS 0.00335f
C2641 VSS.n2070 VSUBS 0.0107f
C2642 VSS.n2071 VSUBS 0.199f
C2643 VSS.n2072 VSUBS 0.0837f
C2644 VSS.n2073 VSUBS 0.0174f
C2645 VSS.t67 VSUBS 0.0109f
C2646 VSS.t108 VSUBS 0.0109f
C2647 VSS.n2074 VSUBS 0.0263f
C2648 VSS.n2075 VSUBS 0.00951f
C2649 VSS.n2076 VSUBS 0.0254f
C2650 VSS.n2077 VSUBS 0.00679f
C2651 VSS.n2078 VSUBS 0.00335f
C2652 VSS.n2079 VSUBS 0.0107f
C2653 VSS.n2080 VSUBS 0.0816f
C2654 VSS.n2081 VSUBS 0.0837f
C2655 VSS.n2082 VSUBS 0.0174f
C2656 VSS.t119 VSUBS 0.0109f
C2657 VSS.t37 VSUBS 0.0109f
C2658 VSS.n2083 VSUBS 0.0263f
C2659 VSS.n2084 VSUBS 0.00951f
C2660 VSS.n2085 VSUBS 0.0254f
C2661 VSS.n2086 VSUBS 0.00679f
C2662 VSS.n2087 VSUBS 0.00335f
C2663 VSS.n2088 VSUBS 0.0107f
C2664 VSS.n2089 VSUBS 0.0816f
C2665 VSS.n2090 VSUBS 0.0837f
C2666 VSS.n2091 VSUBS 0.0174f
C2667 VSS.t47 VSUBS 0.0109f
C2668 VSS.t128 VSUBS 0.0109f
C2669 VSS.n2092 VSUBS 0.0263f
C2670 VSS.n2093 VSUBS 0.00951f
C2671 VSS.n2094 VSUBS 0.0254f
C2672 VSS.n2095 VSUBS 0.00679f
C2673 VSS.n2096 VSUBS 0.00335f
C2674 VSS.n2097 VSUBS 0.0107f
C2675 VSS.n2098 VSUBS 0.0816f
C2676 VSS.n2099 VSUBS 0.0837f
C2677 VSS.n2100 VSUBS 0.0174f
C2678 VSS.t104 VSUBS 0.0109f
C2679 VSS.t24 VSUBS 0.0109f
C2680 VSS.n2101 VSUBS 0.0263f
C2681 VSS.n2102 VSUBS 0.00951f
C2682 VSS.n2103 VSUBS 0.0254f
C2683 VSS.n2104 VSUBS 0.00679f
C2684 VSS.n2105 VSUBS 0.00335f
C2685 VSS.n2106 VSUBS 0.0107f
C2686 VSS.n2107 VSUBS 0.0816f
C2687 VSS.n2108 VSUBS 0.0837f
C2688 VSS.n2109 VSUBS 0.0174f
C2689 VSS.t76 VSUBS 0.0109f
C2690 VSS.t80 VSUBS 0.0109f
C2691 VSS.n2110 VSUBS 0.0263f
C2692 VSS.n2111 VSUBS 0.00951f
C2693 VSS.n2112 VSUBS 0.0254f
C2694 VSS.n2113 VSUBS 0.00679f
C2695 VSS.n2114 VSUBS 0.00335f
C2696 VSS.n2115 VSUBS 0.0107f
C2697 VSS.n2116 VSUBS 0.0816f
C2698 VSS.n2117 VSUBS 0.0837f
C2699 VSS.n2118 VSUBS 0.0174f
C2700 VSS.t41 VSUBS 0.0109f
C2701 VSS.t50 VSUBS 0.0109f
C2702 VSS.n2119 VSUBS 0.0263f
C2703 VSS.n2120 VSUBS 0.00951f
C2704 VSS.n2121 VSUBS 0.0254f
C2705 VSS.n2122 VSUBS 0.00679f
C2706 VSS.n2123 VSUBS 0.00335f
C2707 VSS.n2124 VSUBS 0.0107f
C2708 VSS.n2125 VSUBS 0.0816f
C2709 VSS.n2126 VSUBS 0.0837f
C2710 VSS.n2127 VSUBS 0.0174f
C2711 VSS.t77 VSUBS 0.0109f
C2712 VSS.t71 VSUBS 0.0109f
C2713 VSS.n2128 VSUBS 0.0263f
C2714 VSS.n2129 VSUBS 0.00951f
C2715 VSS.n2130 VSUBS 0.0254f
C2716 VSS.n2131 VSUBS 0.00679f
C2717 VSS.n2132 VSUBS 0.00335f
C2718 VSS.n2133 VSUBS 0.0107f
C2719 VSS.n2134 VSUBS 0.0816f
C2720 VSS.n2135 VSUBS 0.0837f
C2721 VSS.n2136 VSUBS 0.0174f
C2722 VSS.t66 VSUBS 0.0109f
C2723 VSS.t100 VSUBS 0.0109f
C2724 VSS.n2137 VSUBS 0.0263f
C2725 VSS.n2138 VSUBS 0.00951f
C2726 VSS.n2139 VSUBS 0.0254f
C2727 VSS.n2140 VSUBS 0.00679f
C2728 VSS.n2141 VSUBS 0.00335f
C2729 VSS.n2142 VSUBS 0.0107f
C2730 VSS.n2143 VSUBS 0.0816f
C2731 VSS.n2144 VSUBS 0.0837f
C2732 VSS.n2145 VSUBS 0.0174f
C2733 VSS.t94 VSUBS 0.0109f
C2734 VSS.t54 VSUBS 0.0109f
C2735 VSS.n2146 VSUBS 0.0263f
C2736 VSS.n2147 VSUBS 0.00951f
C2737 VSS.n2148 VSUBS 0.0254f
C2738 VSS.n2149 VSUBS 0.00679f
C2739 VSS.n2150 VSUBS 0.00335f
C2740 VSS.n2151 VSUBS 0.0107f
C2741 VSS.n2152 VSUBS 0.0816f
C2742 VSS.n2153 VSUBS 0.0837f
C2743 VSS.n2154 VSUBS 0.0174f
C2744 VSS.t46 VSUBS 0.0109f
C2745 VSS.t126 VSUBS 0.0109f
C2746 VSS.n2155 VSUBS 0.0263f
C2747 VSS.n2156 VSUBS 0.00951f
C2748 VSS.n2157 VSUBS 0.0254f
C2749 VSS.n2158 VSUBS 0.00679f
C2750 VSS.n2159 VSUBS 0.00335f
C2751 VSS.n2160 VSUBS 0.0107f
C2752 VSS.n2161 VSUBS 0.0816f
C2753 VSS.n2162 VSUBS 0.0837f
C2754 VSS.n2163 VSUBS 0.0174f
C2755 VSS.t45 VSUBS 0.0109f
C2756 VSS.t34 VSUBS 0.0109f
C2757 VSS.n2164 VSUBS 0.0263f
C2758 VSS.n2165 VSUBS 0.00951f
C2759 VSS.n2166 VSUBS 0.0254f
C2760 VSS.n2167 VSUBS 0.00679f
C2761 VSS.n2168 VSUBS 0.00335f
C2762 VSS.n2169 VSUBS 0.0107f
C2763 VSS.n2170 VSUBS 0.0816f
C2764 VSS.n2171 VSUBS 0.0837f
C2765 VSS.n2172 VSUBS 0.0174f
C2766 VSS.t116 VSUBS 0.0109f
C2767 VSS.t105 VSUBS 0.0109f
C2768 VSS.n2173 VSUBS 0.0263f
C2769 VSS.n2174 VSUBS 0.00951f
C2770 VSS.n2175 VSUBS 0.0254f
C2771 VSS.n2176 VSUBS 0.00679f
C2772 VSS.n2177 VSUBS 0.00335f
C2773 VSS.n2178 VSUBS 0.0107f
C2774 VSS.n2179 VSUBS 0.0816f
C2775 VSS.n2180 VSUBS 0.0837f
C2776 VSS.n2181 VSUBS 0.0174f
C2777 VSS.t64 VSUBS 0.0109f
C2778 VSS.t31 VSUBS 0.0109f
C2779 VSS.n2182 VSUBS 0.0263f
C2780 VSS.n2183 VSUBS 0.00951f
C2781 VSS.n2184 VSUBS 0.0254f
C2782 VSS.n2185 VSUBS 0.00679f
C2783 VSS.n2186 VSUBS 0.00335f
C2784 VSS.n2187 VSUBS 0.0107f
C2785 VSS.n2188 VSUBS 0.0816f
C2786 VSS.n2189 VSUBS 0.0837f
C2787 VSS.n2190 VSUBS 0.0174f
C2788 VSS.t113 VSUBS 0.0109f
C2789 VSS.t69 VSUBS 0.0109f
C2790 VSS.n2191 VSUBS 0.0263f
C2791 VSS.n2192 VSUBS 0.00951f
C2792 VSS.n2193 VSUBS 0.0254f
C2793 VSS.n2194 VSUBS 0.00679f
C2794 VSS.n2195 VSUBS 0.00335f
C2795 VSS.n2196 VSUBS 0.0107f
C2796 VSS.n2197 VSUBS 0.0816f
C2797 VSS.n2198 VSUBS 0.0837f
C2798 VSS.n2199 VSUBS 0.0174f
C2799 VSS.t61 VSUBS 0.0109f
C2800 VSS.t134 VSUBS 0.0109f
C2801 VSS.n2200 VSUBS 0.0263f
C2802 VSS.n2201 VSUBS 0.00951f
C2803 VSS.n2202 VSUBS 0.0254f
C2804 VSS.n2203 VSUBS 0.00679f
C2805 VSS.n2204 VSUBS 0.00335f
C2806 VSS.n2205 VSUBS 0.0107f
C2807 VSS.n2206 VSUBS 0.0816f
C2808 VSS.n2207 VSUBS 0.0837f
C2809 VSS.n2208 VSUBS 0.0174f
C2810 VSS.t90 VSUBS 0.0109f
C2811 VSS.t68 VSUBS 0.0109f
C2812 VSS.n2209 VSUBS 0.0263f
C2813 VSS.n2210 VSUBS 0.00951f
C2814 VSS.n2211 VSUBS 0.0254f
C2815 VSS.n2212 VSUBS 0.00679f
C2816 VSS.n2213 VSUBS 0.00335f
C2817 VSS.n2214 VSUBS 0.0107f
C2818 VSS.n2215 VSUBS 0.0816f
C2819 VSS.n2216 VSUBS 0.0837f
C2820 VSS.n2217 VSUBS 0.0174f
C2821 VSS.t137 VSUBS 0.0109f
C2822 VSS.t133 VSUBS 0.0109f
C2823 VSS.n2218 VSUBS 0.0263f
C2824 VSS.n2219 VSUBS 0.00951f
C2825 VSS.n2220 VSUBS 0.0254f
C2826 VSS.n2221 VSUBS 0.00679f
C2827 VSS.n2222 VSUBS 0.00335f
C2828 VSS.n2223 VSUBS 0.0107f
C2829 VSS.n2224 VSUBS 0.0816f
C2830 VSS.n2225 VSUBS 0.0837f
C2831 VSS.n2226 VSUBS 0.0174f
C2832 VSS.t79 VSUBS 0.0109f
C2833 VSS.t49 VSUBS 0.0109f
C2834 VSS.n2227 VSUBS 0.0263f
C2835 VSS.n2228 VSUBS 0.00951f
C2836 VSS.n2229 VSUBS 0.0254f
C2837 VSS.n2230 VSUBS 0.00679f
C2838 VSS.n2231 VSUBS 0.00335f
C2839 VSS.n2232 VSUBS 0.0107f
C2840 VSS.n2233 VSUBS 0.0816f
C2841 VSS.n2234 VSUBS 0.0837f
C2842 VSS.n2235 VSUBS 0.0174f
C2843 VSS.t125 VSUBS 0.0109f
C2844 VSS.t121 VSUBS 0.0109f
C2845 VSS.n2236 VSUBS 0.0263f
C2846 VSS.n2237 VSUBS 0.00951f
C2847 VSS.n2238 VSUBS 0.0254f
C2848 VSS.n2239 VSUBS 0.00679f
C2849 VSS.n2240 VSUBS 0.00335f
C2850 VSS.n2241 VSUBS 0.0107f
C2851 VSS.n2242 VSUBS 0.0782f
C2852 VSS.n2244 VSUBS 0.0148f
C2853 VSS.n2245 VSUBS 0.0145f
C2854 VSS.n2246 VSUBS 0.0148f
C2855 VSS.n2247 VSUBS 0.00689f
C2856 VSS.n2248 VSUBS 0.0148f
C2857 VSS.n2249 VSUBS 0.00689f
C2858 VSS.n2250 VSUBS 0.0148f
C2859 VSS.n2251 VSUBS 0.00689f
C2860 VSS.n2252 VSUBS 0.0148f
C2861 VSS.n2253 VSUBS 0.00689f
C2862 VSS.n2254 VSUBS 0.0148f
C2863 VSS.n2255 VSUBS 0.00689f
C2864 VSS.n2256 VSUBS 0.0148f
C2865 VSS.n2257 VSUBS 0.00689f
C2866 VSS.n2258 VSUBS 0.0148f
C2867 VSS.n2259 VSUBS 0.00689f
C2868 VSS.n2260 VSUBS 0.0148f
C2869 VSS.n2261 VSUBS 0.00689f
C2870 VSS.n2262 VSUBS 0.0293f
C2871 VSS.n2263 VSUBS 0.00785f
C2872 VSS.n2264 VSUBS 0.0283f
C2873 VSS.n2265 VSUBS 0.00853f
C2874 VSS.n2266 VSUBS 0.00626f
C2875 VSS.n2267 VSUBS 0.0148f
C2876 VSS.n2268 VSUBS 0.0654f
C2877 VSS.n2269 VSUBS 0.0495f
C2878 VSS.n2270 VSUBS 0.00867f
C2879 VSS.n2271 VSUBS 0.0768f
C2880 VSS.n2272 VSUBS 0.0195f
C2881 VSS.n2273 VSUBS 0.142f
C2882 VSS.n2274 VSUBS 0.114f
C2883 VSS.n2275 VSUBS 0.0235f
C2884 VSS.n2276 VSUBS 0.164f
C2885 VSS.n2277 VSUBS 0.0148f
C2886 VSS.n2278 VSUBS 0.0214f
C2887 VSS.n2280 VSUBS 0.0193f
C2888 VSS.n2281 VSUBS 0.0121f
C2889 VSS.n2283 VSUBS 0.0148f
C2890 VSS.n2284 VSUBS 0.02f
C2891 VSS.n2285 VSUBS 0.0148f
C2892 VSS.n2286 VSUBS 0.0421f
C2893 VSS.n2287 VSUBS 0.00867f
C2894 VSS.n2288 VSUBS 0.0135f
C2895 VSS.n2289 VSUBS 0.0148f
C2896 VSS.n2290 VSUBS 0.0186f
C2897 VSS.n2291 VSUBS 0.0148f
C2898 VSS.n2292 VSUBS 0.0421f
C2899 VSS.n2294 VSUBS 0.00867f
C2900 VSS.n2295 VSUBS 0.0148f
C2901 VSS.n2297 VSUBS 0.0148f
C2902 VSS.n2298 VSUBS 0.0173f
C2903 VSS.n2299 VSUBS 0.0148f
C2904 VSS.n2300 VSUBS 0.0421f
C2905 VSS.n2301 VSUBS 0.00867f
C2906 VSS.n2302 VSUBS 0.0162f
C2907 VSS.n2303 VSUBS 0.0148f
C2908 VSS.n2304 VSUBS 0.0159f
C2909 VSS.n2305 VSUBS 0.0148f
C2910 VSS.n2306 VSUBS 0.0421f
C2911 VSS.n2308 VSUBS 0.00867f
C2912 VSS.n2309 VSUBS 0.0176f
C2913 VSS.n2311 VSUBS 0.0148f
C2914 VSS.n2312 VSUBS 0.0145f
C2915 VSS.n2313 VSUBS 0.0148f
C2916 VSS.n2314 VSUBS 0.0421f
C2917 VSS.n2315 VSUBS 0.00867f
C2918 VSS.n2316 VSUBS 0.019f
C2919 VSS.n2317 VSUBS 0.0148f
C2920 VSS.n2318 VSUBS 0.0131f
C2921 VSS.n2319 VSUBS 0.0148f
C2922 VSS.n2320 VSUBS 0.0421f
C2923 VSS.n2321 VSUBS 0.00867f
C2924 VSS.n2322 VSUBS 0.0204f
C2925 VSS.n2324 VSUBS 0.00867f
C2926 VSS.n2325 VSUBS 0.0217f
C2927 VSS.n2327 VSUBS 0.0148f
C2928 VSS.n2328 VSUBS 0.0117f
C2929 VSS.n2329 VSUBS 0.0148f
C2930 VSS.n2330 VSUBS 0.0421f
C2931 VSS.n2331 VSUBS 0.00867f
C2932 VSS.n2332 VSUBS 0.0231f
C2933 VSS.n2333 VSUBS 0.0148f
C2934 VSS.n2334 VSUBS 0.0104f
C2935 VSS.n2335 VSUBS 0.0148f
C2936 VSS.n2336 VSUBS 0.0421f
C2937 VSS.n2338 VSUBS 0.00867f
C2938 VSS.n2339 VSUBS 0.0235f
C2939 VSS.n2341 VSUBS 0.0148f
C2940 VSS.n2342 VSUBS 0.00897f
C2941 VSS.n2343 VSUBS 0.0148f
C2942 VSS.n2344 VSUBS 0.0421f
C2943 VSS.n2346 VSUBS 0.0148f
C2944 VSS.n2347 VSUBS 0.0159f
C2945 VSS.n2348 VSUBS 0.00867f
C2946 VSS.n2349 VSUBS 0.0224f
C2947 VSS.n2350 VSUBS 0.00863f
C2948 VSS.n2351 VSUBS 0.0421f
C2949 VSS.n2352 VSUBS 0.0148f
C2950 VSS.n2353 VSUBS 0.0173f
C2951 VSS.n2355 VSUBS 0.00867f
C2952 VSS.n2356 VSUBS 0.021f
C2953 VSS.n2357 VSUBS 0.00863f
C2954 VSS.n2358 VSUBS 0.0421f
C2955 VSS.n2360 VSUBS 0.0148f
C2956 VSS.n2361 VSUBS 0.0186f
C2957 VSS.n2362 VSUBS 0.00867f
C2958 VSS.n2363 VSUBS 0.0197f
C2959 VSS.n2364 VSUBS 0.00863f
C2960 VSS.n2365 VSUBS 0.0421f
C2961 VSS.n2366 VSUBS 0.0148f
C2962 VSS.n2367 VSUBS 0.02f
C2963 VSS.n2369 VSUBS 0.00867f
C2964 VSS.n2370 VSUBS 0.0183f
C2965 VSS.n2371 VSUBS 0.00863f
C2966 VSS.n2372 VSUBS 0.0421f
C2967 VSS.n2374 VSUBS 0.0148f
C2968 VSS.n2375 VSUBS 0.0214f
C2969 VSS.n2376 VSUBS 0.00867f
C2970 VSS.n2377 VSUBS 0.0169f
C2971 VSS.n2378 VSUBS 0.00863f
C2972 VSS.n2379 VSUBS 0.0421f
C2973 VSS.n2380 VSUBS 0.0148f
C2974 VSS.n2381 VSUBS 0.0228f
C2975 VSS.n2383 VSUBS 0.00867f
C2976 VSS.n2384 VSUBS 0.0155f
C2977 VSS.n2385 VSUBS 0.00863f
C2978 VSS.n2386 VSUBS 0.0414f
C2979 VSS.n2388 VSUBS 0.0148f
C2980 VSS.n2389 VSUBS 0.0235f
C2981 VSS.n2391 VSUBS 0.00867f
C2982 VSS.n2392 VSUBS 0.00932f
C2983 VSS.n2393 VSUBS 0.0148f
C2984 VSS.n2394 VSUBS 0.206f
C2985 VSS.n2395 VSUBS 0.0148f
C2986 VSS.n2396 VSUBS 0.0228f
C2987 VSS.n2397 VSUBS 0.00867f
C2988 VSS.n2398 VSUBS 0.0107f
C2989 VSS.n2399 VSUBS 0.0148f
C2990 VSS.n2400 VSUBS 0.344f
C2991 VSS.n2401 VSUBS 0.0148f
C2992 VSS.n2402 VSUBS 0.0214f
C2993 VSS.n2404 VSUBS 0.00867f
C2994 VSS.n2405 VSUBS 0.0121f
C2995 VSS.n2407 VSUBS 0.0148f
C2996 VSS.n2408 VSUBS 0.02f
C2997 VSS.n2409 VSUBS 0.0148f
C2998 VSS.n2410 VSUBS 0.397f
C2999 VSS.n2411 VSUBS 0.00867f
C3000 VSS.n2412 VSUBS 0.0135f
C3001 VSS.n2413 VSUBS 0.0148f
C3002 VSS.n2414 VSUBS 0.0186f
C3003 VSS.n2415 VSUBS 0.0148f
C3004 VSS.n2416 VSUBS 0.0603f
C3005 VSS.n2418 VSUBS 0.00867f
C3006 VSS.n2419 VSUBS 0.0148f
C3007 VSS.n2421 VSUBS 0.0148f
C3008 VSS.n2422 VSUBS 0.0173f
C3009 VSS.n2423 VSUBS 0.0148f
C3010 VSS.n2424 VSUBS 0.0421f
C3011 VSS.n2425 VSUBS 0.00867f
C3012 VSS.n2426 VSUBS 0.0162f
C3013 VSS.n2427 VSUBS 0.0148f
C3014 VSS.n2428 VSUBS 0.0159f
C3015 VSS.n2429 VSUBS 0.0148f
C3016 VSS.n2430 VSUBS 0.0421f
C3017 VSS.n2432 VSUBS 0.00867f
C3018 VSS.n2433 VSUBS 0.0176f
C3019 VSS.n2435 VSUBS 0.0148f
C3020 VSS.n2436 VSUBS 0.0145f
C3021 VSS.n2437 VSUBS 0.0148f
C3022 VSS.n2438 VSUBS 0.0421f
C3023 VSS.n2439 VSUBS 0.00867f
C3024 VSS.n2440 VSUBS 0.019f
C3025 VSS.n2441 VSUBS 0.0148f
C3026 VSS.n2442 VSUBS 0.0131f
C3027 VSS.n2443 VSUBS 0.0148f
C3028 VSS.n2444 VSUBS 0.0421f
C3029 VSS.n2445 VSUBS 0.00867f
C3030 VSS.n2446 VSUBS 0.0204f
C3031 VSS.n2448 VSUBS 0.00867f
C3032 VSS.n2449 VSUBS 0.0217f
C3033 VSS.n2451 VSUBS 0.0148f
C3034 VSS.n2452 VSUBS 0.0117f
C3035 VSS.n2453 VSUBS 0.0148f
C3036 VSS.n2454 VSUBS 0.0421f
C3037 VSS.n2455 VSUBS 0.00867f
C3038 VSS.n2456 VSUBS 0.0231f
C3039 VSS.n2457 VSUBS 0.0148f
C3040 VSS.n2458 VSUBS 0.0104f
C3041 VSS.n2459 VSUBS 0.0148f
C3042 VSS.n2460 VSUBS 0.0421f
C3043 VSS.n2462 VSUBS 0.00867f
C3044 VSS.n2463 VSUBS 0.0235f
C3045 VSS.n2465 VSUBS 0.0148f
C3046 VSS.n2466 VSUBS 0.00897f
C3047 VSS.n2467 VSUBS 0.0148f
C3048 VSS.n2468 VSUBS 0.0421f
C3049 VSS.n2470 VSUBS 0.0148f
C3050 VSS.n2471 VSUBS 0.0159f
C3051 VSS.n2472 VSUBS 0.00867f
C3052 VSS.n2473 VSUBS 0.0224f
C3053 VSS.n2474 VSUBS 0.00863f
C3054 VSS.n2475 VSUBS 0.123f
C3055 VSS.n2476 VSUBS 0.0148f
C3056 VSS.n2477 VSUBS 0.0173f
C3057 VSS.n2479 VSUBS 0.00867f
C3058 VSS.n2480 VSUBS 0.021f
C3059 VSS.n2481 VSUBS 0.00863f
C3060 VSS.n2482 VSUBS 0.393f
C3061 VSS.n2484 VSUBS 0.0148f
C3062 VSS.n2485 VSUBS 0.0186f
C3063 VSS.n2486 VSUBS 0.00867f
C3064 VSS.n2487 VSUBS 0.0197f
C3065 VSS.n2488 VSUBS 0.00863f
C3066 VSS.n2489 VSUBS 0.406f
C3067 VSS.n2490 VSUBS 0.0148f
C3068 VSS.n2491 VSUBS 0.02f
C3069 VSS.n2493 VSUBS 0.00867f
C3070 VSS.n2494 VSUBS 0.0183f
C3071 VSS.n2495 VSUBS 0.00863f
C3072 VSS.n2496 VSUBS 0.0845f
C3073 VSS.n2498 VSUBS 0.0148f
C3074 VSS.n2499 VSUBS 0.0214f
C3075 VSS.n2500 VSUBS 0.00867f
C3076 VSS.n2501 VSUBS 0.0169f
C3077 VSS.n2502 VSUBS 0.00863f
C3078 VSS.n2503 VSUBS 0.0421f
C3079 VSS.n2504 VSUBS 0.0148f
C3080 VSS.n2505 VSUBS 0.0228f
C3081 VSS.n2507 VSUBS 0.00867f
C3082 VSS.n2508 VSUBS 0.0155f
C3083 VSS.n2509 VSUBS 0.00863f
C3084 VSS.n2510 VSUBS 0.0421f
C3085 VSS.n2512 VSUBS 0.0148f
C3086 VSS.n2513 VSUBS 0.0235f
C3087 VSS.n2515 VSUBS 0.00867f
C3088 VSS.n2516 VSUBS 0.00932f
C3089 VSS.n2517 VSUBS 0.0148f
C3090 VSS.n2518 VSUBS 0.0421f
C3091 VSS.n2519 VSUBS 0.0148f
C3092 VSS.n2520 VSUBS 0.0228f
C3093 VSS.n2521 VSUBS 0.00867f
C3094 VSS.n2522 VSUBS 0.0107f
C3095 VSS.n2523 VSUBS 0.0148f
C3096 VSS.n2524 VSUBS 0.0421f
C3097 VSS.n2525 VSUBS 0.0148f
C3098 VSS.n2526 VSUBS 0.0214f
C3099 VSS.n2528 VSUBS 0.00867f
C3100 VSS.n2529 VSUBS 0.0121f
C3101 VSS.n2531 VSUBS 0.0148f
C3102 VSS.n2532 VSUBS 0.02f
C3103 VSS.n2533 VSUBS 0.0148f
C3104 VSS.n2534 VSUBS 0.0421f
C3105 VSS.n2535 VSUBS 0.00867f
C3106 VSS.n2536 VSUBS 0.0135f
C3107 VSS.n2537 VSUBS 0.0148f
C3108 VSS.n2538 VSUBS 0.0186f
C3109 VSS.n2539 VSUBS 0.0148f
C3110 VSS.n2540 VSUBS 0.0421f
C3111 VSS.n2542 VSUBS 0.00867f
C3112 VSS.n2543 VSUBS 0.0148f
C3113 VSS.n2545 VSUBS 0.0148f
C3114 VSS.n2546 VSUBS 0.0173f
C3115 VSS.n2547 VSUBS 0.0148f
C3116 VSS.n2548 VSUBS 0.0421f
C3117 VSS.n2549 VSUBS 0.00867f
C3118 VSS.n2550 VSUBS 0.0162f
C3119 VSS.n2551 VSUBS 0.0148f
C3120 VSS.n2552 VSUBS 0.0159f
C3121 VSS.n2553 VSUBS 0.0148f
C3122 VSS.n2554 VSUBS 0.0766f
C3123 VSS.n2556 VSUBS 0.00867f
C3124 VSS.n2557 VSUBS 0.0176f
C3125 VSS.n2559 VSUBS 0.0148f
C3126 VSS.n2560 VSUBS 0.0145f
C3127 VSS.n2561 VSUBS 0.0148f
C3128 VSS.n2562 VSUBS 0.406f
C3129 VSS.n2563 VSUBS 0.00867f
C3130 VSS.n2564 VSUBS 0.019f
C3131 VSS.n2565 VSUBS 0.0148f
C3132 VSS.n2566 VSUBS 0.0131f
C3133 VSS.n2567 VSUBS 0.0148f
C3134 VSS.n2568 VSUBS 0.38f
C3135 VSS.n2570 VSUBS 0.00867f
C3136 VSS.n2571 VSUBS 0.0204f
C3137 VSS.n2572 VSUBS 0.00867f
C3138 VSS.n2573 VSUBS 0.0217f
C3139 VSS.n2575 VSUBS 0.0148f
C3140 VSS.n2576 VSUBS 0.0117f
C3141 VSS.n2577 VSUBS 0.0148f
C3142 VSS.n2578 VSUBS 0.144f
C3143 VSS.n2579 VSUBS 0.00867f
C3144 VSS.n2580 VSUBS 0.0231f
C3145 VSS.n2581 VSUBS 0.0148f
C3146 VSS.n2582 VSUBS 0.0104f
C3147 VSS.n2583 VSUBS 0.0148f
C3148 VSS.n2584 VSUBS 0.0421f
C3149 VSS.n2586 VSUBS 0.00867f
C3150 VSS.n2587 VSUBS 0.0235f
C3151 VSS.n2589 VSUBS 0.0148f
C3152 VSS.n2590 VSUBS 0.00897f
C3153 VSS.n2591 VSUBS 0.0148f
C3154 VSS.n2592 VSUBS 0.0421f
C3155 VSS.n2594 VSUBS 0.0148f
C3156 VSS.n2595 VSUBS 0.0159f
C3157 VSS.n2596 VSUBS 0.00867f
C3158 VSS.n2597 VSUBS 0.0224f
C3159 VSS.n2598 VSUBS 0.00863f
C3160 VSS.n2599 VSUBS 0.0421f
C3161 VSS.n2600 VSUBS 0.0148f
C3162 VSS.n2601 VSUBS 0.0173f
C3163 VSS.n2603 VSUBS 0.00867f
C3164 VSS.n2604 VSUBS 0.021f
C3165 VSS.n2605 VSUBS 0.00863f
C3166 VSS.n2606 VSUBS 0.0421f
C3167 VSS.n2608 VSUBS 0.0148f
C3168 VSS.n2609 VSUBS 0.0186f
C3169 VSS.n2610 VSUBS 0.00867f
C3170 VSS.n2611 VSUBS 0.0197f
C3171 VSS.n2612 VSUBS 0.00863f
C3172 VSS.n2613 VSUBS 0.0421f
C3173 VSS.n2614 VSUBS 0.0148f
C3174 VSS.n2615 VSUBS 0.02f
C3175 VSS.n2617 VSUBS 0.00867f
C3176 VSS.n2618 VSUBS 0.0183f
C3177 VSS.n2619 VSUBS 0.00863f
C3178 VSS.n2620 VSUBS 0.0421f
C3179 VSS.n2622 VSUBS 0.0148f
C3180 VSS.n2623 VSUBS 0.0214f
C3181 VSS.n2624 VSUBS 0.00867f
C3182 VSS.n2625 VSUBS 0.0169f
C3183 VSS.n2626 VSUBS 0.00863f
C3184 VSS.n2627 VSUBS 0.0421f
C3185 VSS.n2628 VSUBS 0.0148f
C3186 VSS.n2629 VSUBS 0.0228f
C3187 VSS.n2631 VSUBS 0.00867f
C3188 VSS.n2632 VSUBS 0.0155f
C3189 VSS.n2633 VSUBS 0.00863f
C3190 VSS.n2634 VSUBS 0.0565f
C3191 VSS.n2636 VSUBS 0.0148f
C3192 VSS.n2637 VSUBS 0.0235f
C3193 VSS.n2639 VSUBS 0.00867f
C3194 VSS.n2640 VSUBS 0.00932f
C3195 VSS.n2641 VSUBS 0.0148f
C3196 VSS.n2642 VSUBS 0.392f
C3197 VSS.n2643 VSUBS 0.0148f
C3198 VSS.n2644 VSUBS 0.0228f
C3199 VSS.n2645 VSUBS 0.00867f
C3200 VSS.n2646 VSUBS 0.0107f
C3201 VSS.n2647 VSUBS 0.0148f
C3202 VSS.n2648 VSUBS 0.344f
C3203 VSS.n2649 VSUBS 0.0148f
C3204 VSS.n2650 VSUBS 0.0214f
C3205 VSS.n2652 VSUBS 0.00867f
C3206 VSS.n2653 VSUBS 0.0121f
C3207 VSS.n2655 VSUBS 0.0148f
C3208 VSS.n2656 VSUBS 0.02f
C3209 VSS.n2657 VSUBS 0.0148f
C3210 VSS.n2658 VSUBS 0.215f
C3211 VSS.n2659 VSUBS 0.00867f
C3212 VSS.n2660 VSUBS 0.0135f
C3213 VSS.n2661 VSUBS 0.0148f
C3214 VSS.n2662 VSUBS 0.0186f
C3215 VSS.n2663 VSUBS 0.0148f
C3216 VSS.n2664 VSUBS 0.0409f
C3217 VSS.n2666 VSUBS 0.00867f
C3218 VSS.n2667 VSUBS 0.0148f
C3219 VSS.n2669 VSUBS 0.0148f
C3220 VSS.n2670 VSUBS 0.0173f
C3221 VSS.n2671 VSUBS 0.0148f
C3222 VSS.n2672 VSUBS 0.0421f
C3223 VSS.n2673 VSUBS 0.00867f
C3224 VSS.n2674 VSUBS 0.0162f
C3225 VSS.n2675 VSUBS 0.0148f
C3226 VSS.n2676 VSUBS 0.0159f
C3227 VSS.n2677 VSUBS 0.0148f
C3228 VSS.n2678 VSUBS 0.0421f
C3229 VSS.n2680 VSUBS 0.00867f
C3230 VSS.n2681 VSUBS 0.0176f
C3231 VSS.n2683 VSUBS 0.0148f
C3232 VSS.n2684 VSUBS 0.0145f
C3233 VSS.n2685 VSUBS 0.0148f
C3234 VSS.n2686 VSUBS 0.0421f
C3235 VSS.n2687 VSUBS 0.00867f
C3236 VSS.n2688 VSUBS 0.019f
C3237 VSS.n2689 VSUBS 0.0148f
C3238 VSS.n2690 VSUBS 0.0131f
C3239 VSS.n2691 VSUBS 0.0148f
C3240 VSS.n2692 VSUBS 0.0421f
C3241 VSS.n2694 VSUBS 0.00867f
C3242 VSS.n2695 VSUBS 0.0204f
C3243 VSS.n2696 VSUBS 0.00867f
C3244 VSS.n2697 VSUBS 0.0217f
C3245 VSS.n2699 VSUBS 0.0148f
C3246 VSS.n2700 VSUBS 0.0117f
C3247 VSS.n2701 VSUBS 0.0148f
C3248 VSS.n2702 VSUBS 0.0421f
C3249 VSS.n2703 VSUBS 0.00867f
C3250 VSS.n2704 VSUBS 0.0231f
C3251 VSS.n2705 VSUBS 0.0148f
C3252 VSS.n2706 VSUBS 0.0104f
C3253 VSS.n2707 VSUBS 0.0148f
C3254 VSS.n2708 VSUBS 0.0421f
C3255 VSS.n2710 VSUBS 0.00867f
C3256 VSS.n2711 VSUBS 0.0235f
C3257 VSS.n2713 VSUBS 0.0148f
C3258 VSS.n2714 VSUBS 0.00897f
C3259 VSS.n2715 VSUBS 0.0148f
C3260 VSS.n2716 VSUBS 0.0466f
C3261 VSS.n2718 VSUBS 0.0148f
C3262 VSS.n2719 VSUBS 0.0159f
C3263 VSS.n2720 VSUBS 0.00867f
C3264 VSS.n2721 VSUBS 0.0224f
C3265 VSS.n2722 VSUBS 0.00863f
C3266 VSS.n2723 VSUBS 0.369f
C3267 VSS.n2724 VSUBS 0.0148f
C3268 VSS.n2725 VSUBS 0.0173f
C3269 VSS.n2727 VSUBS 0.00867f
C3270 VSS.n2728 VSUBS 0.021f
C3271 VSS.n2729 VSUBS 0.00863f
C3272 VSS.n2730 VSUBS 0.344f
C3273 VSS.n2732 VSUBS 0.0148f
C3274 VSS.n2733 VSUBS 0.0186f
C3275 VSS.n2734 VSUBS 0.00867f
C3276 VSS.n2735 VSUBS 0.0197f
C3277 VSS.n2736 VSUBS 0.00863f
C3278 VSS.n2737 VSUBS 0.25f
C3279 VSS.n2738 VSUBS 0.0148f
C3280 VSS.n2739 VSUBS 0.02f
C3281 VSS.n2741 VSUBS 0.00867f
C3282 VSS.n2742 VSUBS 0.0183f
C3283 VSS.n2743 VSUBS 0.00863f
C3284 VSS.n2744 VSUBS 0.0396f
C3285 VSS.n2746 VSUBS 0.0148f
C3286 VSS.n2747 VSUBS 0.0214f
C3287 VSS.n2748 VSUBS 0.00867f
C3288 VSS.n2749 VSUBS 0.0169f
C3289 VSS.n2750 VSUBS 0.00863f
C3290 VSS.n2751 VSUBS 0.0421f
C3291 VSS.n2752 VSUBS 0.0148f
C3292 VSS.n2753 VSUBS 0.0228f
C3293 VSS.n2755 VSUBS 0.00867f
C3294 VSS.n2756 VSUBS 0.0155f
C3295 VSS.n2757 VSUBS 0.00863f
C3296 VSS.n2758 VSUBS 0.0421f
C3297 VSS.n2760 VSUBS 0.0148f
C3298 VSS.n2761 VSUBS 0.0235f
C3299 VSS.n2763 VSUBS 0.00867f
C3300 VSS.n2764 VSUBS 0.00932f
C3301 VSS.n2765 VSUBS 0.0148f
C3302 VSS.n2766 VSUBS 0.0421f
C3303 VSS.n2767 VSUBS 0.0148f
C3304 VSS.n2768 VSUBS 0.0228f
C3305 VSS.n2769 VSUBS 0.00867f
C3306 VSS.n2770 VSUBS 0.0107f
C3307 VSS.n2771 VSUBS 0.0148f
C3308 VSS.n2772 VSUBS 0.0421f
C3309 VSS.n2773 VSUBS 0.0148f
C3310 VSS.n2774 VSUBS 0.0214f
C3311 VSS.n2776 VSUBS 0.00867f
C3312 VSS.n2777 VSUBS 0.0121f
C3313 VSS.n2779 VSUBS 0.0148f
C3314 VSS.n2780 VSUBS 0.02f
C3315 VSS.n2781 VSUBS 0.0148f
C3316 VSS.n2782 VSUBS 0.0421f
C3317 VSS.n2783 VSUBS 0.00867f
C3318 VSS.n2784 VSUBS 0.0135f
C3319 VSS.n2785 VSUBS 0.0148f
C3320 VSS.n2786 VSUBS 0.0186f
C3321 VSS.n2787 VSUBS 0.0148f
C3322 VSS.n2788 VSUBS 0.0421f
C3323 VSS.n2790 VSUBS 0.00867f
C3324 VSS.n2791 VSUBS 0.0148f
C3325 VSS.n2793 VSUBS 0.0148f
C3326 VSS.n2794 VSUBS 0.0173f
C3327 VSS.n2795 VSUBS 0.0148f
C3328 VSS.n2796 VSUBS 0.0417f
C3329 VSS.n2797 VSUBS 0.00867f
C3330 VSS.n2798 VSUBS 0.0162f
C3331 VSS.n2799 VSUBS 0.0148f
C3332 VSS.n2800 VSUBS 0.0159f
C3333 VSS.n2801 VSUBS 0.0148f
C3334 VSS.n2802 VSUBS 0.34f
C3335 VSS.n2804 VSUBS 0.00867f
C3336 VSS.n2805 VSUBS 0.0176f
C3337 VSS.n2807 VSUBS 0.0148f
C3338 VSS.n2808 VSUBS 0.0145f
C3339 VSS.n2809 VSUBS 0.0148f
C3340 VSS.n2810 VSUBS 0.344f
C3341 VSS.n2811 VSUBS 0.00867f
C3342 VSS.n2812 VSUBS 0.019f
C3343 VSS.n2813 VSUBS 0.0148f
C3344 VSS.n2814 VSUBS 0.0131f
C3345 VSS.n2815 VSUBS 0.0148f
C3346 VSS.n2816 VSUBS 0.284f
C3347 VSS.n2818 VSUBS 0.00867f
C3348 VSS.n2819 VSUBS 0.0204f
C3349 VSS.n2820 VSUBS 0.00867f
C3350 VSS.n2821 VSUBS 0.0217f
C3351 VSS.n2823 VSUBS 0.0148f
C3352 VSS.n2824 VSUBS 0.0117f
C3353 VSS.n2825 VSUBS 0.0148f
C3354 VSS.n2826 VSUBS 0.0391f
C3355 VSS.n2827 VSUBS 0.00867f
C3356 VSS.n2828 VSUBS 0.0231f
C3357 VSS.n2829 VSUBS 0.0148f
C3358 VSS.n2830 VSUBS 0.0104f
C3359 VSS.n2831 VSUBS 0.0148f
C3360 VSS.n2832 VSUBS 0.0421f
C3361 VSS.n2834 VSUBS 0.00867f
C3362 VSS.n2835 VSUBS 0.0235f
C3363 VSS.n2837 VSUBS 0.0148f
C3364 VSS.n2838 VSUBS 0.00897f
C3365 VSS.n2839 VSUBS 0.0148f
C3366 VSS.n2840 VSUBS 0.0421f
C3367 VSS.n2842 VSUBS 0.0148f
C3368 VSS.n2843 VSUBS 0.0159f
C3369 VSS.n2844 VSUBS 0.00867f
C3370 VSS.n2845 VSUBS 0.0224f
C3371 VSS.n2846 VSUBS 0.00863f
C3372 VSS.n2847 VSUBS 0.0421f
C3373 VSS.n2848 VSUBS 0.0148f
C3374 VSS.n2849 VSUBS 0.0173f
C3375 VSS.n2851 VSUBS 0.00867f
C3376 VSS.n2852 VSUBS 0.021f
C3377 VSS.n2853 VSUBS 0.00863f
C3378 VSS.n2854 VSUBS 0.0421f
C3379 VSS.n2856 VSUBS 0.0148f
C3380 VSS.n2857 VSUBS 0.0186f
C3381 VSS.n2858 VSUBS 0.00867f
C3382 VSS.n2859 VSUBS 0.0197f
C3383 VSS.n2860 VSUBS 0.00863f
C3384 VSS.n2861 VSUBS 0.0421f
C3385 VSS.n2862 VSUBS 0.0148f
C3386 VSS.n2863 VSUBS 0.02f
C3387 VSS.n2865 VSUBS 0.00867f
C3388 VSS.n2866 VSUBS 0.0183f
C3389 VSS.n2867 VSUBS 0.00863f
C3390 VSS.n2868 VSUBS 0.0421f
C3391 VSS.n2870 VSUBS 0.0148f
C3392 VSS.n2871 VSUBS 0.0214f
C3393 VSS.n2872 VSUBS 0.0193f
C3394 VSS.n2873 VSUBS 0.0169f
C3395 VSS.n2874 VSUBS 0.00863f
C3396 VSS.n2875 VSUBS 0.0421f
C3397 VSS.n2876 VSUBS 0.0148f
C3398 VSS.n2877 VSUBS 0.0228f
C3399 VSS.n2878 VSUBS 0.021f
C3400 VSS.n2879 VSUBS 0.0612f
C3401 VSS.n2880 VSUBS 0.0148f
C3402 VSS.n2881 VSUBS 0.00842f
C3403 VSS.n2882 VSUBS 0.0148f
C3404 VSS.n2883 VSUBS 0.00842f
C3405 VSS.n2884 VSUBS 0.0148f
C3406 VSS.n2885 VSUBS 0.00842f
C3407 VSS.n2886 VSUBS 0.0148f
C3408 VSS.n2887 VSUBS 0.00842f
C3409 VSS.n2888 VSUBS 0.0148f
C3410 VSS.n2889 VSUBS 0.00842f
C3411 VSS.n2890 VSUBS 0.0148f
C3412 VSS.n2891 VSUBS 0.00842f
C3413 VSS.n2892 VSUBS 0.0148f
C3414 VSS.n2893 VSUBS 0.00842f
C3415 VSS.n2894 VSUBS 0.0148f
C3416 VSS.n2895 VSUBS 0.00842f
C3417 VSS.n2896 VSUBS 0.0293f
C3418 VSS.n2897 VSUBS 0.00963f
C3419 VSS.n2898 VSUBS 0.0148f
C3420 VSS.n2899 VSUBS 1.72f
C3421 VSS.n2900 VSUBS 1.72f
C3422 VSS.n2901 VSUBS 1.72f
C3423 VSS.n2902 VSUBS 1.72f
C3424 VSS.n2903 VSUBS 1.72f
C3425 VSS.n2904 VSUBS 0.985f
C3426 VSS.t23 VSUBS 0.859f
C3427 VSS.n2905 VSUBS 1.59f
C3428 VSS.n2906 VSUBS 1.72f
C3429 VSS.n2907 VSUBS 2.11f
C3430 VSS.t0 VSUBS 0.859f
C3431 VSS.n2908 VSUBS 1.87f
C3432 VSS.n2909 VSUBS 3.35f
C3433 VSS.n2910 VSUBS 3.14f
C3434 VSS.n2911 VSUBS 0.0074f
C3435 VSS.n2912 VSUBS 0.0074f
C3436 VSS.n2913 VSUBS 0.0283f
C3437 VSS.n2914 VSUBS 0.0587f
C3438 VSS.n2915 VSUBS 0.055f
C3439 VSS.n2916 VSUBS 0.0405f
C3440 VSS.n2917 VSUBS 0.216f
C3441 VSS.n2918 VSUBS 0.0694f
C3442 VSS.n2919 VSUBS 0.0709f
C3443 VSS.n2920 VSUBS 0.00867f
C3444 VSS.n2921 VSUBS 0.0474f
C3445 VSS.n2922 VSUBS 0.0389f
C3446 VSS.n2923 VSUBS 0.00867f
C3447 VSS.n2924 VSUBS 0.0406f
C3448 VSS.n2925 VSUBS 0.0384f
C3449 VSS.n2926 VSUBS 0.0625f
C3450 VSS.n2927 VSUBS 0.00867f
C3451 VSS.n2928 VSUBS 0.0406f
C3452 VSS.n2929 VSUBS 0.0384f
C3453 VSS.n2930 VSUBS 0.0302f
C3454 VSS.n2931 VSUBS 0.00867f
C3455 VSS.n2932 VSUBS 0.0406f
C3456 VSS.n2933 VSUBS 0.0384f
C3457 VSS.n2934 VSUBS 0.0302f
C3458 VSS.n2935 VSUBS 0.00867f
C3459 VSS.n2936 VSUBS 0.0406f
C3460 VSS.n2937 VSUBS 0.0384f
C3461 VSS.n2938 VSUBS 0.0302f
C3462 VSS.n2939 VSUBS 0.00867f
C3463 VSS.n2940 VSUBS 0.0214f
C3464 VSS.n2941 VSUBS 0.0426f
C3465 VSS.n2942 VSUBS 0.00867f
C3466 VSS.n2943 VSUBS 0.0406f
C3467 VSS.n2944 VSUBS 0.0373f
C3468 VSS.n2945 VSUBS 0.0302f
C3469 VSS.n2946 VSUBS 0.00867f
C3470 VSS.n2947 VSUBS 0.0406f
C3471 VSS.n2948 VSUBS 0.0384f
C3472 VSS.n2949 VSUBS 0.0302f
C3473 VSS.n2950 VSUBS 0.00867f
C3474 VSS.n2951 VSUBS 0.0406f
C3475 VSS.n2952 VSUBS 0.0384f
C3476 VSS.n2953 VSUBS 0.0302f
C3477 VSS.n2954 VSUBS 0.00867f
C3478 VSS.n2955 VSUBS 0.0406f
C3479 VSS.n2956 VSUBS 0.0384f
C3480 VSS.n2957 VSUBS 0.0302f
C3481 VSS.n2958 VSUBS 0.00867f
C3482 VSS.n2959 VSUBS 0.0406f
C3483 VSS.n2960 VSUBS 0.0384f
C3484 VSS.n2961 VSUBS 0.0302f
C3485 VSS.n2962 VSUBS 0.00867f
C3486 VSS.n2963 VSUBS 0.0406f
C3487 VSS.n2964 VSUBS 0.0384f
C3488 VSS.n2965 VSUBS 0.0302f
C3489 VSS.n2966 VSUBS 0.00867f
C3490 VSS.n2967 VSUBS 0.0406f
C3491 VSS.n2968 VSUBS 0.0384f
C3492 VSS.n2969 VSUBS 0.0302f
C3493 VSS.n2970 VSUBS 0.0195f
C3494 VSS.n2971 VSUBS 0.0406f
C3495 VSS.n2972 VSUBS 0.0384f
C3496 VSS.n2973 VSUBS 0.0302f
C3497 VSS.n2974 VSUBS 0.079f
C3498 VSS.n2975 VSUBS 0.0302f
C3499 VSS.n2976 VSUBS 0.0548f
C3500 VSS.n2977 VSUBS 0.0508f
C3501 VSS.n2978 VSUBS 0.0728f
C3502 VSS.n2979 VSUBS 0.0529f
C3503 VSS.n2980 VSUBS 0.0234f
C3504 VSS.n2981 VSUBS 0.0321f
C3505 VSS.n2983 VSUBS 0.0193f
C3506 VSS.n2984 VSUBS 0.0162f
C3507 VSS.n2985 VSUBS 0.0153f
C3508 VSS.n2986 VSUBS 0.024f
C3509 VSS.n2987 VSUBS 0.00867f
C3510 VSS.n2988 VSUBS 0.0162f
C3511 VSS.n2989 VSUBS 0.0153f
C3512 VSS.n2990 VSUBS 0.024f
C3513 VSS.n2992 VSUBS 0.00867f
C3514 VSS.n2993 VSUBS 0.0162f
C3515 VSS.n2994 VSUBS 0.0153f
C3516 VSS.n2995 VSUBS 0.024f
C3517 VSS.n2997 VSUBS 0.00867f
C3518 VSS.n2998 VSUBS 0.0162f
C3519 VSS.n2999 VSUBS 0.0153f
C3520 VSS.n3000 VSUBS 0.024f
C3521 VSS.n3001 VSUBS 0.00867f
C3522 VSS.n3002 VSUBS 0.0162f
C3523 VSS.n3003 VSUBS 0.0153f
C3524 VSS.n3004 VSUBS 0.024f
C3525 VSS.n3006 VSUBS 0.00867f
C3526 VSS.n3007 VSUBS 0.0162f
C3527 VSS.n3008 VSUBS 0.0153f
C3528 VSS.n3009 VSUBS 0.024f
C3529 VSS.n3010 VSUBS 0.00867f
C3530 VSS.n3011 VSUBS 0.0162f
C3531 VSS.n3012 VSUBS 0.00867f
C3532 VSS.n3013 VSUBS 0.0162f
C3533 VSS.n3014 VSUBS 0.0153f
C3534 VSS.n3015 VSUBS 0.024f
C3535 VSS.n3017 VSUBS 0.00867f
C3536 VSS.n3018 VSUBS 0.0162f
C3537 VSS.n3019 VSUBS 0.0153f
C3538 VSS.n3020 VSUBS 0.024f
C3539 VSS.n3021 VSUBS 0.00867f
C3540 VSS.n3022 VSUBS 0.0162f
C3541 VSS.n3023 VSUBS 0.0153f
C3542 VSS.n3024 VSUBS 0.024f
C3543 VSS.n3026 VSUBS 0.00867f
C3544 VSS.n3027 VSUBS 0.0162f
C3545 VSS.n3028 VSUBS 0.0153f
C3546 VSS.n3029 VSUBS 0.0275f
C3547 VSS.n3030 VSUBS 0.00867f
C3548 VSS.n3031 VSUBS 0.0162f
C3549 VSS.n3032 VSUBS 0.0153f
C3550 VSS.n3033 VSUBS 0.348f
C3551 VSS.n3035 VSUBS 0.00867f
C3552 VSS.n3036 VSUBS 0.0162f
C3553 VSS.n3037 VSUBS 0.0153f
C3554 VSS.n3038 VSUBS 0.319f
C3555 VSS.n3039 VSUBS 0.00867f
C3556 VSS.n3040 VSUBS 0.0162f
C3557 VSS.n3041 VSUBS 0.0153f
C3558 VSS.n3042 VSUBS 0.222f
C3559 VSS.n3044 VSUBS 0.00867f
C3560 VSS.n3045 VSUBS 0.0162f
C3561 VSS.n3046 VSUBS 0.0153f
C3562 VSS.n3047 VSUBS 0.0226f
C3563 VSS.n3049 VSUBS 0.00867f
C3564 VSS.n3050 VSUBS 0.0155f
C3565 VSS.n3051 VSUBS 0.0153f
C3566 VSS.n3052 VSUBS 0.024f
C3567 VSS.n3053 VSUBS 0.00867f
C3568 VSS.n3054 VSUBS 0.016f
C3569 VSS.n3055 VSUBS 0.0153f
C3570 VSS.n3056 VSUBS 0.024f
C3571 VSS.n3058 VSUBS 0.00867f
C3572 VSS.n3059 VSUBS 0.0162f
C3573 VSS.n3060 VSUBS 0.0153f
C3574 VSS.n3061 VSUBS 0.024f
C3575 VSS.n3062 VSUBS 0.00867f
C3576 VSS.n3063 VSUBS 0.0162f
C3577 VSS.n3064 VSUBS 0.0153f
C3578 VSS.n3065 VSUBS 0.024f
C3579 VSS.n3067 VSUBS 0.00867f
C3580 VSS.n3068 VSUBS 0.0162f
C3581 VSS.n3069 VSUBS 0.0153f
C3582 VSS.n3070 VSUBS 0.024f
C3583 VSS.n3071 VSUBS 0.00867f
C3584 VSS.n3072 VSUBS 0.0162f
C3585 VSS.n3073 VSUBS 0.0153f
C3586 VSS.n3074 VSUBS 0.024f
C3587 VSS.n3076 VSUBS 0.00867f
C3588 VSS.n3077 VSUBS 0.0162f
C3589 VSS.n3078 VSUBS 0.0153f
C3590 VSS.n3079 VSUBS 0.024f
C3591 VSS.n3080 VSUBS 0.00867f
C3592 VSS.n3081 VSUBS 0.0162f
C3593 VSS.n3082 VSUBS 0.0153f
C3594 VSS.n3083 VSUBS 0.319f
C3595 VSS.n3085 VSUBS 0.00867f
C3596 VSS.n3086 VSUBS 0.0162f
C3597 VSS.n3087 VSUBS 0.0153f
C3598 VSS.n3088 VSUBS 0.319f
C3599 VSS.n3089 VSUBS 0.00867f
C3600 VSS.n3090 VSUBS 0.0162f
C3601 VSS.n3091 VSUBS 0.00867f
C3602 VSS.n3092 VSUBS 0.0162f
C3603 VSS.n3093 VSUBS 0.0153f
C3604 VSS.n3094 VSUBS 0.255f
C3605 VSS.n3096 VSUBS 0.00867f
C3606 VSS.n3097 VSUBS 0.0162f
C3607 VSS.n3098 VSUBS 0.0153f
C3608 VSS.n3099 VSUBS 0.0222f
C3609 VSS.n3100 VSUBS 0.00867f
C3610 VSS.n3101 VSUBS 0.0162f
C3611 VSS.n3102 VSUBS 0.0153f
C3612 VSS.n3103 VSUBS 0.024f
C3613 VSS.n3105 VSUBS 0.00867f
C3614 VSS.n3106 VSUBS 0.0162f
C3615 VSS.n3107 VSUBS 0.0153f
C3616 VSS.n3108 VSUBS 0.024f
C3617 VSS.n3109 VSUBS 0.00867f
C3618 VSS.n3110 VSUBS 0.0162f
C3619 VSS.n3111 VSUBS 0.0153f
C3620 VSS.n3112 VSUBS 0.024f
C3621 VSS.n3114 VSUBS 0.00867f
C3622 VSS.n3115 VSUBS 0.0162f
C3623 VSS.n3116 VSUBS 0.0153f
C3624 VSS.n3117 VSUBS 0.024f
C3625 VSS.n3118 VSUBS 0.00867f
C3626 VSS.n3119 VSUBS 0.0162f
C3627 VSS.n3120 VSUBS 0.0153f
C3628 VSS.n3121 VSUBS 0.024f
C3629 VSS.n3123 VSUBS 0.00867f
C3630 VSS.n3124 VSUBS 0.0162f
C3631 VSS.n3125 VSUBS 0.0153f
C3632 VSS.n3126 VSUBS 0.024f
C3633 VSS.n3128 VSUBS 0.00867f
C3634 VSS.n3129 VSUBS 0.0155f
C3635 VSS.n3130 VSUBS 0.0153f
C3636 VSS.n3131 VSUBS 0.0225f
C3637 VSS.n3132 VSUBS 0.00867f
C3638 VSS.n3133 VSUBS 0.016f
C3639 VSS.n3134 VSUBS 0.0153f
C3640 VSS.n3135 VSUBS 0.287f
C3641 VSS.n3137 VSUBS 0.00867f
C3642 VSS.n3138 VSUBS 0.0162f
C3643 VSS.n3139 VSUBS 0.0153f
C3644 VSS.n3140 VSUBS 0.319f
C3645 VSS.n3141 VSUBS 0.00867f
C3646 VSS.n3142 VSUBS 0.0162f
C3647 VSS.n3143 VSUBS 0.0153f
C3648 VSS.n3144 VSUBS 0.287f
C3649 VSS.n3146 VSUBS 0.00867f
C3650 VSS.n3147 VSUBS 0.0162f
C3651 VSS.n3148 VSUBS 0.0153f
C3652 VSS.n3149 VSUBS 0.0225f
C3653 VSS.n3150 VSUBS 0.00867f
C3654 VSS.n3151 VSUBS 0.0162f
C3655 VSS.n3152 VSUBS 0.0153f
C3656 VSS.n3153 VSUBS 0.024f
C3657 VSS.n3155 VSUBS 0.00867f
C3658 VSS.n3156 VSUBS 0.0162f
C3659 VSS.n3157 VSUBS 0.0153f
C3660 VSS.n3158 VSUBS 0.024f
C3661 VSS.n3159 VSUBS 0.00867f
C3662 VSS.n3160 VSUBS 0.0162f
C3663 VSS.n3161 VSUBS 0.0153f
C3664 VSS.n3162 VSUBS 0.024f
C3665 VSS.n3164 VSUBS 0.00867f
C3666 VSS.n3165 VSUBS 0.0162f
C3667 VSS.n3166 VSUBS 0.0153f
C3668 VSS.n3167 VSUBS 0.024f
C3669 VSS.n3168 VSUBS 0.00867f
C3670 VSS.n3169 VSUBS 0.0162f
C3671 VSS.n3170 VSUBS 0.00867f
C3672 VSS.n3171 VSUBS 0.0162f
C3673 VSS.n3172 VSUBS 0.0153f
C3674 VSS.n3173 VSUBS 0.024f
C3675 VSS.n3175 VSUBS 0.00867f
C3676 VSS.n3176 VSUBS 0.0162f
C3677 VSS.n3177 VSUBS 0.0153f
C3678 VSS.n3178 VSUBS 0.024f
C3679 VSS.n3179 VSUBS 0.00867f
C3680 VSS.n3180 VSUBS 0.0162f
C3681 VSS.n3181 VSUBS 0.0153f
C3682 VSS.n3182 VSUBS 0.0222f
C3683 VSS.n3184 VSUBS 0.00867f
C3684 VSS.n3185 VSUBS 0.0162f
C3685 VSS.n3186 VSUBS 0.0153f
C3686 VSS.n3187 VSUBS 0.255f
C3687 VSS.n3188 VSUBS 0.00867f
C3688 VSS.n3189 VSUBS 0.0162f
C3689 VSS.n3190 VSUBS 0.0153f
C3690 VSS.n3191 VSUBS 0.319f
C3691 VSS.n3193 VSUBS 0.00867f
C3692 VSS.n3194 VSUBS 0.0162f
C3693 VSS.n3195 VSUBS 0.0153f
C3694 VSS.n3196 VSUBS 0.319f
C3695 VSS.n3197 VSUBS 0.00867f
C3696 VSS.n3198 VSUBS 0.0162f
C3697 VSS.n3199 VSUBS 0.0153f
C3698 VSS.n3200 VSUBS 0.024f
C3699 VSS.n3202 VSUBS 0.00867f
C3700 VSS.n3203 VSUBS 0.0162f
C3701 VSS.n3204 VSUBS 0.0153f
C3702 VSS.n3205 VSUBS 0.024f
C3703 VSS.n3207 VSUBS 0.00867f
C3704 VSS.n3208 VSUBS 0.0155f
C3705 VSS.n3209 VSUBS 0.0153f
C3706 VSS.n3210 VSUBS 0.024f
C3707 VSS.n3211 VSUBS 0.00867f
C3708 VSS.n3212 VSUBS 0.016f
C3709 VSS.n3213 VSUBS 0.0153f
C3710 VSS.n3214 VSUBS 0.024f
C3711 VSS.n3216 VSUBS 0.00867f
C3712 VSS.n3217 VSUBS 0.0162f
C3713 VSS.n3218 VSUBS 0.0153f
C3714 VSS.n3219 VSUBS 0.024f
C3715 VSS.n3220 VSUBS 0.00867f
C3716 VSS.n3221 VSUBS 0.0162f
C3717 VSS.n3222 VSUBS 0.0153f
C3718 VSS.n3223 VSUBS 0.024f
C3719 VSS.n3225 VSUBS 0.00867f
C3720 VSS.n3226 VSUBS 0.0162f
C3721 VSS.n3227 VSUBS 0.0153f
C3722 VSS.n3228 VSUBS 0.024f
C3723 VSS.n3229 VSUBS 0.00867f
C3724 VSS.n3230 VSUBS 0.0162f
C3725 VSS.n3231 VSUBS 0.0153f
C3726 VSS.n3232 VSUBS 0.0226f
C3727 VSS.n3234 VSUBS 0.00867f
C3728 VSS.n3235 VSUBS 0.0162f
C3729 VSS.n3236 VSUBS 0.0153f
C3730 VSS.n3237 VSUBS 0.222f
C3731 VSS.n3238 VSUBS 0.00867f
C3732 VSS.n3239 VSUBS 0.0162f
C3733 VSS.n3240 VSUBS 0.0153f
C3734 VSS.n3241 VSUBS 0.319f
C3735 VSS.n3243 VSUBS 0.00867f
C3736 VSS.n3244 VSUBS 0.0162f
C3737 VSS.n3245 VSUBS 0.0153f
C3738 VSS.n3246 VSUBS 0.348f
C3739 VSS.n3247 VSUBS 0.00867f
C3740 VSS.n3248 VSUBS 0.0162f
C3741 VSS.n3249 VSUBS 0.00867f
C3742 VSS.n3250 VSUBS 0.0162f
C3743 VSS.n3251 VSUBS 0.0153f
C3744 VSS.n3252 VSUBS 0.0275f
C3745 VSS.n3254 VSUBS 0.00867f
C3746 VSS.n3255 VSUBS 0.0162f
C3747 VSS.n3256 VSUBS 0.0153f
C3748 VSS.n3257 VSUBS 0.024f
C3749 VSS.n3258 VSUBS 0.00867f
C3750 VSS.n3259 VSUBS 0.0162f
C3751 VSS.n3260 VSUBS 0.0153f
C3752 VSS.n3261 VSUBS 0.024f
C3753 VSS.n3263 VSUBS 0.00867f
C3754 VSS.n3264 VSUBS 0.0162f
C3755 VSS.n3265 VSUBS 0.0153f
C3756 VSS.n3266 VSUBS 0.024f
C3757 VSS.n3267 VSUBS 0.00867f
C3758 VSS.n3268 VSUBS 0.0162f
C3759 VSS.n3269 VSUBS 0.0153f
C3760 VSS.n3270 VSUBS 0.024f
C3761 VSS.n3272 VSUBS 0.00867f
C3762 VSS.n3273 VSUBS 0.0162f
C3763 VSS.n3274 VSUBS 0.0153f
C3764 VSS.n3275 VSUBS 0.024f
C3765 VSS.n3276 VSUBS 0.00867f
C3766 VSS.n3277 VSUBS 0.0162f
C3767 VSS.n3278 VSUBS 0.0153f
C3768 VSS.n3279 VSUBS 0.024f
C3769 VSS.n3281 VSUBS 0.00867f
C3770 VSS.n3282 VSUBS 0.0162f
C3771 VSS.n3283 VSUBS 0.0153f
C3772 VSS.n3284 VSUBS 0.0235f
C3773 VSS.n3286 VSUBS 0.00867f
C3774 VSS.n3287 VSUBS 0.0155f
C3775 VSS.n3288 VSUBS 0.0153f
C3776 VSS.n3289 VSUBS 0.188f
C3777 VSS.n3290 VSUBS 0.00867f
C3778 VSS.n3291 VSUBS 0.016f
C3779 VSS.n3292 VSUBS 0.0153f
C3780 VSS.n3293 VSUBS 0.319f
C3781 VSS.n3295 VSUBS 0.00867f
C3782 VSS.n3296 VSUBS 0.0162f
C3783 VSS.n3297 VSUBS 0.0153f
C3784 VSS.n3298 VSUBS 0.373f
C3785 VSS.n3299 VSUBS 0.00867f
C3786 VSS.n3300 VSUBS 0.0162f
C3787 VSS.n3301 VSUBS 0.0153f
C3788 VSS.n3302 VSUBS 0.0348f
C3789 VSS.n3304 VSUBS 0.00867f
C3790 VSS.n3305 VSUBS 0.0162f
C3791 VSS.n3306 VSUBS 0.0153f
C3792 VSS.n3307 VSUBS 0.024f
C3793 VSS.n3308 VSUBS 0.00867f
C3794 VSS.n3309 VSUBS 0.0162f
C3795 VSS.n3310 VSUBS 0.0153f
C3796 VSS.n3311 VSUBS 0.024f
C3797 VSS.n3313 VSUBS 0.00867f
C3798 VSS.n3314 VSUBS 0.0162f
C3799 VSS.n3315 VSUBS 0.0153f
C3800 VSS.n3316 VSUBS 0.024f
C3801 VSS.n3317 VSUBS 0.00867f
C3802 VSS.n3318 VSUBS 0.0162f
C3803 VSS.n3319 VSUBS 0.0153f
C3804 VSS.n3320 VSUBS 0.024f
C3805 VSS.n3322 VSUBS 0.00867f
C3806 VSS.n3323 VSUBS 0.0162f
C3807 VSS.n3324 VSUBS 0.0153f
C3808 VSS.n3325 VSUBS 0.024f
C3809 VSS.n3326 VSUBS 0.00867f
C3810 VSS.n3327 VSUBS 0.0162f
C3811 VSS.n3328 VSUBS 0.00867f
C3812 VSS.n3329 VSUBS 0.0162f
C3813 VSS.n3330 VSUBS 0.0153f
C3814 VSS.n3331 VSUBS 0.024f
C3815 VSS.n3333 VSUBS 0.00867f
C3816 VSS.n3334 VSUBS 0.0162f
C3817 VSS.n3335 VSUBS 0.0153f
C3818 VSS.n3336 VSUBS 0.024f
C3819 VSS.n3337 VSUBS 0.00867f
C3820 VSS.n3338 VSUBS 0.0162f
C3821 VSS.n3339 VSUBS 0.0153f
C3822 VSS.n3340 VSUBS 0.024f
C3823 VSS.n3342 VSUBS 0.00867f
C3824 VSS.n3343 VSUBS 0.0162f
C3825 VSS.n3344 VSUBS 0.0153f
C3826 VSS.n3345 VSUBS 0.024f
C3827 VSS.n3346 VSUBS 0.00867f
C3828 VSS.n3347 VSUBS 0.0162f
C3829 VSS.n3348 VSUBS 0.0153f
C3830 VSS.n3349 VSUBS 0.024f
C3831 VSS.n3351 VSUBS 0.00867f
C3832 VSS.n3352 VSUBS 0.0162f
C3833 VSS.n3353 VSUBS 0.0153f
C3834 VSS.n3354 VSUBS 0.024f
C3835 VSS.n3355 VSUBS 0.00867f
C3836 VSS.n3356 VSUBS 0.0162f
C3837 VSS.n3357 VSUBS 0.0153f
C3838 VSS.n3358 VSUBS 0.024f
C3839 VSS.t2 VSUBS 0.859f
C3840 VSS.n3359 VSUBS 1.87f
C3841 VSS.n3360 VSUBS 3.55f
C3842 VSS.n3362 VSUBS 0.0193f
C3843 VSS.n3363 VSUBS 0.0162f
C3844 VSS.n3364 VSUBS 0.0153f
C3845 VSS.n3365 VSUBS 0.024f
C3846 VSS.n3366 VSUBS 0.0234f
C3847 VSS.n3367 VSUBS 0.024f
C3848 VSS.n3368 VSUBS 0.0868f
C3849 VSS.n3369 VSUBS 0.0534f
C3850 VSS.n3370 VSUBS 0.0636f
C3851 VSS.n3371 VSUBS 0.0572f
C3852 VSS.n3372 VSUBS 0.0195f
C3853 VSS.n3373 VSUBS 0.0347f
C3854 VSS.n3374 VSUBS 0.0472f
C3855 VSS.n3375 VSUBS 0.0354f
C3856 VSS.n3376 VSUBS 1.3f
C3857 VSS.n3377 VSUBS 0.00867f
C3858 VSS.n3378 VSUBS 0.0347f
C3859 VSS.n3379 VSUBS 0.0328f
C3860 VSS.n3380 VSUBS 0.0354f
C3861 VSS.n3381 VSUBS 1.72f
C3862 VSS.n3382 VSUBS 0.00867f
C3863 VSS.n3383 VSUBS 0.0347f
C3864 VSS.n3384 VSUBS 0.0328f
C3865 VSS.n3385 VSUBS 0.0354f
C3866 VSS.n3386 VSUBS 1.72f
C3867 VSS.n3387 VSUBS 0.00867f
C3868 VSS.n3388 VSUBS 0.0347f
C3869 VSS.n3389 VSUBS 0.0328f
C3870 VSS.n3390 VSUBS 0.0354f
C3871 VSS.n3391 VSUBS 1.72f
C3872 VSS.n3392 VSUBS 0.00867f
C3873 VSS.n3393 VSUBS 0.0347f
C3874 VSS.n3394 VSUBS 0.0328f
C3875 VSS.n3395 VSUBS 0.0354f
C3876 VSS.t10 VSUBS 0.859f
C3877 VSS.n3396 VSUBS 0.998f
C3878 VSS.n3397 VSUBS 0.00867f
C3879 VSS.n3398 VSUBS 0.0347f
C3880 VSS.n3399 VSUBS 0.0328f
C3881 VSS.n3400 VSUBS 0.0354f
C3882 VSS.n3401 VSUBS 1.58f
C3883 VSS.n3402 VSUBS 0.00867f
C3884 VSS.n3403 VSUBS 0.0337f
C3885 VSS.n3404 VSUBS 0.0328f
C3886 VSS.n3405 VSUBS 0.0354f
C3887 VSS.n3406 VSUBS 1.72f
C3888 VSS.n3407 VSUBS 0.00867f
C3889 VSS.n3408 VSUBS 0.0337f
C3890 VSS.n3409 VSUBS 0.0328f
C3891 VSS.n3410 VSUBS 0.0354f
C3892 VSS.n3411 VSUBS 1.72f
C3893 VSS.n3412 VSUBS 0.00867f
C3894 VSS.n3413 VSUBS 0.0347f
C3895 VSS.n3414 VSUBS 0.0328f
C3896 VSS.n3415 VSUBS 0.0354f
C3897 VSS.n3416 VSUBS 1.58f
C3898 VSS.n3417 VSUBS 0.00867f
C3899 VSS.n3418 VSUBS 0.0347f
C3900 VSS.n3419 VSUBS 0.0328f
C3901 VSS.n3420 VSUBS 0.0354f
C3902 VSS.t14 VSUBS 0.859f
C3903 VSS.n3421 VSUBS 0.998f
C3904 VSS.n3422 VSUBS 0.00867f
C3905 VSS.n3423 VSUBS 0.0347f
C3906 VSS.n3424 VSUBS 0.0328f
C3907 VSS.n3425 VSUBS 0.0354f
C3908 VSS.n3426 VSUBS 1.72f
C3909 VSS.n3427 VSUBS 0.00867f
C3910 VSS.n3428 VSUBS 0.0347f
C3911 VSS.n3429 VSUBS 0.0328f
C3912 VSS.n3430 VSUBS 0.0354f
C3913 VSS.n3431 VSUBS 1.72f
C3914 VSS.n3432 VSUBS 0.00867f
C3915 VSS.n3433 VSUBS 0.0347f
C3916 VSS.n3434 VSUBS 0.0328f
C3917 VSS.n3435 VSUBS 0.0354f
C3918 VSS.n3436 VSUBS 1.72f
C3919 VSS.n3437 VSUBS 0.00867f
C3920 VSS.n3438 VSUBS 0.0347f
C3921 VSS.n3439 VSUBS 0.0328f
C3922 VSS.n3440 VSUBS 0.0589f
C3923 VSS.n3441 VSUBS 1.3f
C3924 VSS.n3442 VSUBS 0.00867f
C3925 VSS.n3443 VSUBS 0.0347f
C3926 VSS.n3444 VSUBS 0.0328f
C3927 VSS.n3445 VSUBS 0.114f
C3928 VSS.n3446 VSUBS 0.0195f
C3929 VSS.n3447 VSUBS 0.0347f
C3930 VSS.n3448 VSUBS 0.0511f
C3931 VSS.n3449 VSUBS 0.0903f
C3932 VSS.n3450 VSUBS 0.435f
C3933 VSS.n3451 VSUBS 0.466f
C3934 VSS.n3452 VSUBS 0.487f
C3935 VSS.n3453 VSUBS 0.511f
C3936 VSS.n3454 VSUBS 0.452f
C3937 ndrv.n0 VSUBS 0.899f
C3938 ndrv.n1 VSUBS 1.26f
C3939 ndrv.n2 VSUBS 1.26f
C3940 ndrv.n3 VSUBS 1.26f
C3941 ndrv.n4 VSUBS 1.26f
C3942 ndrv.n5 VSUBS 1.26f
C3943 ndrv.n6 VSUBS 1.26f
C3944 ndrv.n7 VSUBS 1.26f
C3945 ndrv.n8 VSUBS 1.26f
C3946 ndrv.n9 VSUBS 2.92f
C3947 ndrv.n10 VSUBS 1.26f
C3948 ndrv.n11 VSUBS 1.26f
C3949 ndrv.n12 VSUBS 1.26f
C3950 ndrv.n13 VSUBS 1.26f
C3951 ndrv.n14 VSUBS 1.26f
C3952 ndrv.n15 VSUBS 1.26f
C3953 ndrv.n16 VSUBS 1.26f
C3954 ndrv.n17 VSUBS 1.26f
C3955 ndrv.n18 VSUBS 1.26f
C3956 ndrv.n19 VSUBS 0.66f
C3957 ndrv.n20 VSUBS 6.69f
C3958 ndrv.n21 VSUBS 5.64f
C3959 ndrv.n22 VSUBS 0.63f
C3960 ndrv.n23 VSUBS 3.01f
C3961 ndrv.t22 VSUBS 0.152f
C3962 ndrv.t13 VSUBS 0.152f
C3963 ndrv.t70 VSUBS 0.152f
C3964 ndrv.t29 VSUBS 0.152f
C3965 ndrv.t18 VSUBS 0.152f
C3966 ndrv.t100 VSUBS 0.152f
C3967 ndrv.t90 VSUBS 0.152f
C3968 ndrv.t9 VSUBS 0.152f
C3969 ndrv.t33 VSUBS 0.152f
C3970 ndrv.t113 VSUBS 0.152f
C3971 ndrv.t61 VSUBS 0.152f
C3972 ndrv.t57 VSUBS 0.152f
C3973 ndrv.t96 VSUBS 0.152f
C3974 ndrv.t87 VSUBS 0.152f
C3975 ndrv.t60 VSUBS 0.152f
C3976 ndrv.t66 VSUBS 0.152f
C3977 ndrv.t71 VSUBS 0.152f
C3978 ndrv.t37 VSUBS 0.152f
C3979 ndrv.t43 VSUBS 0.152f
C3980 ndrv.t83 VSUBS 0.152f
C3981 ndrv.t91 VSUBS 0.152f
C3982 ndrv.t11 VSUBS 0.152f
C3983 ndrv.t92 VSUBS 0.152f
C3984 ndrv.t103 VSUBS 0.152f
C3985 ndrv.t21 VSUBS 0.152f
C3986 ndrv.t32 VSUBS 0.152f
C3987 ndrv.t73 VSUBS 0.152f
C3988 ndrv.t106 VSUBS 0.152f
C3989 ndrv.t24 VSUBS 0.152f
C3990 ndrv.t68 VSUBS 0.152f
C3991 ndrv.t76 VSUBS 0.152f
C3992 ndrv.t3 VSUBS 0.152f
C3993 ndrv.t47 VSUBS 0.152f
C3994 ndrv.t69 VSUBS 0.152f
C3995 ndrv.t0 VSUBS 0.152f
C3996 ndrv.t4 VSUBS 0.152f
C3997 ndrv.t58 VSUBS 0.152f
C3998 ndrv.t88 VSUBS 0.152f
C3999 ndrv.t12 VSUBS 0.152f
C4000 ndrv.t16 VSUBS 0.152f
C4001 ndrv.n24 VSUBS 1.26f
C4002 ndrv.t36 VSUBS 0.152f
C4003 ndrv.t98 VSUBS 0.152f
C4004 ndrv.t26 VSUBS 0.152f
C4005 ndrv.t89 VSUBS 0.152f
C4006 ndrv.t79 VSUBS 0.152f
C4007 ndrv.t25 VSUBS 0.152f
C4008 ndrv.t40 VSUBS 0.152f
C4009 ndrv.t108 VSUBS 0.152f
C4010 ndrv.t34 VSUBS 0.152f
C4011 ndrv.t95 VSUBS 0.152f
C4012 ndrv.t114 VSUBS 0.152f
C4013 ndrv.t53 VSUBS 0.152f
C4014 ndrv.t104 VSUBS 0.152f
C4015 ndrv.t48 VSUBS 0.152f
C4016 ndrv.t15 VSUBS 0.152f
C4017 ndrv.t82 VSUBS 0.152f
C4018 ndrv.t42 VSUBS 0.152f
C4019 ndrv.t110 VSUBS 0.152f
C4020 ndrv.t118 VSUBS 0.152f
C4021 ndrv.t59 VSUBS 0.152f
C4022 ndrv.t65 VSUBS 0.152f
C4023 ndrv.t6 VSUBS 0.152f
C4024 ndrv.t62 VSUBS 0.152f
C4025 ndrv.t1 VSUBS 0.152f
C4026 ndrv.t111 VSUBS 0.152f
C4027 ndrv.t51 VSUBS 0.152f
C4028 ndrv.t99 VSUBS 0.152f
C4029 ndrv.t44 VSUBS 0.152f
C4030 ndrv.t64 VSUBS 0.152f
C4031 ndrv.t5 VSUBS 0.152f
C4032 ndrv.t74 VSUBS 0.152f
C4033 ndrv.t14 VSUBS 0.152f
C4034 ndrv.t80 VSUBS 0.152f
C4035 ndrv.t27 VSUBS 0.152f
C4036 ndrv.t45 VSUBS 0.152f
C4037 ndrv.t112 VSUBS 0.152f
C4038 ndrv.t52 VSUBS 0.152f
C4039 ndrv.t117 VSUBS 0.152f
C4040 ndrv.t93 VSUBS 0.152f
C4041 ndrv.t39 VSUBS 0.152f
C4042 ndrv.t105 VSUBS 0.152f
C4043 ndrv.t49 VSUBS 0.152f
C4044 ndrv.t17 VSUBS 0.152f
C4045 ndrv.t84 VSUBS 0.152f
C4046 ndrv.t107 VSUBS 0.152f
C4047 ndrv.t50 VSUBS 0.152f
C4048 ndrv.t115 VSUBS 0.152f
C4049 ndrv.t54 VSUBS 0.152f
C4050 ndrv.t35 VSUBS 0.152f
C4051 ndrv.t97 VSUBS 0.152f
C4052 ndrv.t41 VSUBS 0.152f
C4053 ndrv.t109 VSUBS 0.152f
C4054 ndrv.t81 VSUBS 0.152f
C4055 ndrv.t28 VSUBS 0.152f
C4056 ndrv.t116 VSUBS 0.152f
C4057 ndrv.t56 VSUBS 0.152f
C4058 ndrv.t38 VSUBS 0.152f
C4059 ndrv.t101 VSUBS 0.152f
C4060 ndrv.t77 VSUBS 0.152f
C4061 ndrv.t19 VSUBS 0.152f
C4062 ndrv.t85 VSUBS 0.152f
C4063 ndrv.t30 VSUBS 0.152f
C4064 ndrv.t8 VSUBS 0.152f
C4065 ndrv.t72 VSUBS 0.152f
C4066 ndrv.t55 VSUBS 0.152f
C4067 ndrv.t119 VSUBS 0.152f
C4068 ndrv.t78 VSUBS 0.152f
C4069 ndrv.t23 VSUBS 0.152f
C4070 ndrv.t7 VSUBS 0.152f
C4071 ndrv.t67 VSUBS 0.152f
C4072 ndrv.t10 VSUBS 0.152f
C4073 ndrv.t63 VSUBS 0.152f
C4074 ndrv.t102 VSUBS 0.152f
C4075 ndrv.t20 VSUBS 0.152f
C4076 ndrv.t31 VSUBS 0.152f
C4077 ndrv.t75 VSUBS 0.171f
C4078 ndrv.t2 VSUBS 0.152f
C4079 ndrv.t46 VSUBS 0.152f
C4080 ndrv.t86 VSUBS 0.152f
C4081 ndrv.t94 VSUBS 0.152f
C4082 VOUT.n0 VSUBS 0.047f
C4083 VOUT.t481 VSUBS 0.0294f
C4084 VOUT.n1 VSUBS 0.1f
C4085 VOUT.n2 VSUBS 0.0264f
C4086 VOUT.n3 VSUBS 0.071f
C4087 VOUT.n4 VSUBS 0.0182f
C4088 VOUT.n5 VSUBS 0.0089f
C4089 VOUT.n6 VSUBS 0.0347f
C4090 VOUT.n7 VSUBS 0.337f
C4091 VOUT.n8 VSUBS 0.047f
C4092 VOUT.t514 VSUBS 0.0294f
C4093 VOUT.t465 VSUBS 0.0294f
C4094 VOUT.n9 VSUBS 0.0711f
C4095 VOUT.n10 VSUBS 0.0264f
C4096 VOUT.n11 VSUBS 0.071f
C4097 VOUT.n12 VSUBS 0.0182f
C4098 VOUT.n13 VSUBS 0.0089f
C4099 VOUT.n14 VSUBS 0.029f
C4100 VOUT.n15 VSUBS 0.22f
C4101 VOUT.n16 VSUBS 0.226f
C4102 VOUT.n17 VSUBS 0.047f
C4103 VOUT.t362 VSUBS 0.0294f
C4104 VOUT.t472 VSUBS 0.0294f
C4105 VOUT.n18 VSUBS 0.0711f
C4106 VOUT.n19 VSUBS 0.0264f
C4107 VOUT.n20 VSUBS 0.071f
C4108 VOUT.n21 VSUBS 0.0182f
C4109 VOUT.n22 VSUBS 0.0089f
C4110 VOUT.n23 VSUBS 0.029f
C4111 VOUT.n24 VSUBS 0.22f
C4112 VOUT.n25 VSUBS 0.226f
C4113 VOUT.n26 VSUBS 0.047f
C4114 VOUT.t459 VSUBS 0.0294f
C4115 VOUT.t387 VSUBS 0.0294f
C4116 VOUT.n27 VSUBS 0.0711f
C4117 VOUT.n28 VSUBS 0.0264f
C4118 VOUT.n29 VSUBS 0.071f
C4119 VOUT.n30 VSUBS 0.0182f
C4120 VOUT.n31 VSUBS 0.0089f
C4121 VOUT.n32 VSUBS 0.029f
C4122 VOUT.n33 VSUBS 0.22f
C4123 VOUT.n34 VSUBS 0.226f
C4124 VOUT.n35 VSUBS 0.047f
C4125 VOUT.t53 VSUBS 0.0294f
C4126 VOUT.t431 VSUBS 0.0294f
C4127 VOUT.n36 VSUBS 0.0711f
C4128 VOUT.n37 VSUBS 0.0264f
C4129 VOUT.n38 VSUBS 0.071f
C4130 VOUT.n39 VSUBS 0.0182f
C4131 VOUT.n40 VSUBS 0.0089f
C4132 VOUT.n41 VSUBS 0.029f
C4133 VOUT.n42 VSUBS 0.22f
C4134 VOUT.n43 VSUBS 0.226f
C4135 VOUT.n44 VSUBS 0.047f
C4136 VOUT.t448 VSUBS 0.0294f
C4137 VOUT.t452 VSUBS 0.0294f
C4138 VOUT.n45 VSUBS 0.0711f
C4139 VOUT.n46 VSUBS 0.0264f
C4140 VOUT.n47 VSUBS 0.071f
C4141 VOUT.n48 VSUBS 0.0182f
C4142 VOUT.n49 VSUBS 0.0089f
C4143 VOUT.n50 VSUBS 0.029f
C4144 VOUT.n51 VSUBS 0.22f
C4145 VOUT.n52 VSUBS 0.226f
C4146 VOUT.n53 VSUBS 0.047f
C4147 VOUT.t84 VSUBS 0.0294f
C4148 VOUT.t354 VSUBS 0.0294f
C4149 VOUT.n54 VSUBS 0.0711f
C4150 VOUT.n55 VSUBS 0.0264f
C4151 VOUT.n56 VSUBS 0.071f
C4152 VOUT.n57 VSUBS 0.0182f
C4153 VOUT.n58 VSUBS 0.0089f
C4154 VOUT.n59 VSUBS 0.029f
C4155 VOUT.n60 VSUBS 0.22f
C4156 VOUT.n61 VSUBS 0.226f
C4157 VOUT.n62 VSUBS 0.047f
C4158 VOUT.t479 VSUBS 0.0294f
C4159 VOUT.t447 VSUBS 0.0294f
C4160 VOUT.n63 VSUBS 0.0711f
C4161 VOUT.n64 VSUBS 0.0264f
C4162 VOUT.n65 VSUBS 0.071f
C4163 VOUT.n66 VSUBS 0.0182f
C4164 VOUT.n67 VSUBS 0.0089f
C4165 VOUT.n68 VSUBS 0.029f
C4166 VOUT.n69 VSUBS 0.22f
C4167 VOUT.n70 VSUBS 0.226f
C4168 VOUT.n71 VSUBS 0.047f
C4169 VOUT.t435 VSUBS 0.0294f
C4170 VOUT.t31 VSUBS 0.0294f
C4171 VOUT.n72 VSUBS 0.0711f
C4172 VOUT.n73 VSUBS 0.0264f
C4173 VOUT.n74 VSUBS 0.071f
C4174 VOUT.n75 VSUBS 0.0182f
C4175 VOUT.n76 VSUBS 0.0089f
C4176 VOUT.n77 VSUBS 0.029f
C4177 VOUT.n78 VSUBS 0.22f
C4178 VOUT.n79 VSUBS 0.226f
C4179 VOUT.n80 VSUBS 0.047f
C4180 VOUT.t89 VSUBS 0.0294f
C4181 VOUT.t35 VSUBS 0.0294f
C4182 VOUT.n81 VSUBS 0.0711f
C4183 VOUT.n82 VSUBS 0.0264f
C4184 VOUT.n83 VSUBS 0.071f
C4185 VOUT.n84 VSUBS 0.0182f
C4186 VOUT.n85 VSUBS 0.0089f
C4187 VOUT.n86 VSUBS 0.029f
C4188 VOUT.n87 VSUBS 0.22f
C4189 VOUT.n88 VSUBS 0.226f
C4190 VOUT.n89 VSUBS 0.047f
C4191 VOUT.t444 VSUBS 0.0294f
C4192 VOUT.t50 VSUBS 0.0294f
C4193 VOUT.n90 VSUBS 0.0711f
C4194 VOUT.n91 VSUBS 0.0264f
C4195 VOUT.n92 VSUBS 0.071f
C4196 VOUT.n93 VSUBS 0.0182f
C4197 VOUT.n94 VSUBS 0.0089f
C4198 VOUT.n95 VSUBS 0.029f
C4199 VOUT.n96 VSUBS 0.22f
C4200 VOUT.n97 VSUBS 0.226f
C4201 VOUT.n98 VSUBS 0.047f
C4202 VOUT.t426 VSUBS 0.0294f
C4203 VOUT.t407 VSUBS 0.0294f
C4204 VOUT.n99 VSUBS 0.0711f
C4205 VOUT.n100 VSUBS 0.0264f
C4206 VOUT.n101 VSUBS 0.071f
C4207 VOUT.n102 VSUBS 0.0182f
C4208 VOUT.n103 VSUBS 0.0089f
C4209 VOUT.n104 VSUBS 0.029f
C4210 VOUT.n105 VSUBS 0.22f
C4211 VOUT.n106 VSUBS 0.226f
C4212 VOUT.n107 VSUBS 0.047f
C4213 VOUT.t477 VSUBS 0.0294f
C4214 VOUT.t484 VSUBS 0.0294f
C4215 VOUT.n108 VSUBS 0.0711f
C4216 VOUT.n109 VSUBS 0.0264f
C4217 VOUT.n110 VSUBS 0.071f
C4218 VOUT.n111 VSUBS 0.0182f
C4219 VOUT.n112 VSUBS 0.0089f
C4220 VOUT.n113 VSUBS 0.029f
C4221 VOUT.n114 VSUBS 0.22f
C4222 VOUT.n115 VSUBS 0.226f
C4223 VOUT.n116 VSUBS 0.047f
C4224 VOUT.t10 VSUBS 0.0294f
C4225 VOUT.t2 VSUBS 0.0294f
C4226 VOUT.n117 VSUBS 0.0711f
C4227 VOUT.n118 VSUBS 0.0264f
C4228 VOUT.n119 VSUBS 0.071f
C4229 VOUT.n120 VSUBS 0.0182f
C4230 VOUT.n121 VSUBS 0.0089f
C4231 VOUT.n122 VSUBS 0.029f
C4232 VOUT.n123 VSUBS 0.22f
C4233 VOUT.n124 VSUBS 0.226f
C4234 VOUT.n125 VSUBS 0.047f
C4235 VOUT.t382 VSUBS 0.0294f
C4236 VOUT.t402 VSUBS 0.0294f
C4237 VOUT.n126 VSUBS 0.0711f
C4238 VOUT.n127 VSUBS 0.0264f
C4239 VOUT.n128 VSUBS 0.071f
C4240 VOUT.n129 VSUBS 0.0182f
C4241 VOUT.n130 VSUBS 0.0089f
C4242 VOUT.n131 VSUBS 0.029f
C4243 VOUT.n132 VSUBS 0.22f
C4244 VOUT.n133 VSUBS 0.226f
C4245 VOUT.n134 VSUBS 0.047f
C4246 VOUT.t108 VSUBS 0.0294f
C4247 VOUT.t383 VSUBS 0.0294f
C4248 VOUT.n135 VSUBS 0.0711f
C4249 VOUT.n136 VSUBS 0.0264f
C4250 VOUT.n137 VSUBS 0.071f
C4251 VOUT.n138 VSUBS 0.0182f
C4252 VOUT.n139 VSUBS 0.0089f
C4253 VOUT.n140 VSUBS 0.029f
C4254 VOUT.n141 VSUBS 0.22f
C4255 VOUT.n142 VSUBS 0.226f
C4256 VOUT.n143 VSUBS 0.047f
C4257 VOUT.t410 VSUBS 0.0294f
C4258 VOUT.t473 VSUBS 0.0294f
C4259 VOUT.n144 VSUBS 0.0711f
C4260 VOUT.n145 VSUBS 0.0264f
C4261 VOUT.n146 VSUBS 0.071f
C4262 VOUT.n147 VSUBS 0.0182f
C4263 VOUT.n148 VSUBS 0.0089f
C4264 VOUT.n149 VSUBS 0.029f
C4265 VOUT.n150 VSUBS 0.22f
C4266 VOUT.n151 VSUBS 0.226f
C4267 VOUT.n152 VSUBS 0.047f
C4268 VOUT.t0 VSUBS 0.0294f
C4269 VOUT.t136 VSUBS 0.0294f
C4270 VOUT.n153 VSUBS 0.0711f
C4271 VOUT.n154 VSUBS 0.0264f
C4272 VOUT.n155 VSUBS 0.071f
C4273 VOUT.n156 VSUBS 0.0182f
C4274 VOUT.n157 VSUBS 0.0089f
C4275 VOUT.n158 VSUBS 0.029f
C4276 VOUT.n159 VSUBS 0.22f
C4277 VOUT.n160 VSUBS 0.226f
C4278 VOUT.n161 VSUBS 0.047f
C4279 VOUT.t30 VSUBS 0.0294f
C4280 VOUT.t424 VSUBS 0.0294f
C4281 VOUT.n162 VSUBS 0.0711f
C4282 VOUT.n163 VSUBS 0.0264f
C4283 VOUT.n164 VSUBS 0.071f
C4284 VOUT.n165 VSUBS 0.0182f
C4285 VOUT.n166 VSUBS 0.0089f
C4286 VOUT.n167 VSUBS 0.029f
C4287 VOUT.n168 VSUBS 0.22f
C4288 VOUT.n169 VSUBS 0.226f
C4289 VOUT.n170 VSUBS 0.047f
C4290 VOUT.t347 VSUBS 0.0294f
C4291 VOUT.t449 VSUBS 0.0294f
C4292 VOUT.n171 VSUBS 0.0711f
C4293 VOUT.n172 VSUBS 0.0264f
C4294 VOUT.n173 VSUBS 0.071f
C4295 VOUT.n174 VSUBS 0.0182f
C4296 VOUT.n175 VSUBS 0.0089f
C4297 VOUT.n176 VSUBS 0.029f
C4298 VOUT.n177 VSUBS 0.22f
C4299 VOUT.n178 VSUBS 0.226f
C4300 VOUT.n179 VSUBS 0.047f
C4301 VOUT.t49 VSUBS 0.0294f
C4302 VOUT.n180 VSUBS 0.1f
C4303 VOUT.n181 VSUBS 0.0264f
C4304 VOUT.n182 VSUBS 0.071f
C4305 VOUT.n183 VSUBS 0.0182f
C4306 VOUT.n184 VSUBS 0.0089f
C4307 VOUT.n185 VSUBS 0.029f
C4308 VOUT.n186 VSUBS 0.22f
C4309 VOUT.n187 VSUBS 0.113f
C4310 VOUT.n188 VSUBS 0.047f
C4311 VOUT.t451 VSUBS 0.0294f
C4312 VOUT.n189 VSUBS 0.1f
C4313 VOUT.n190 VSUBS 0.0264f
C4314 VOUT.n191 VSUBS 0.071f
C4315 VOUT.n192 VSUBS 0.0182f
C4316 VOUT.n193 VSUBS 0.0089f
C4317 VOUT.n194 VSUBS 0.034f
C4318 VOUT.n195 VSUBS 0.322f
C4319 VOUT.n196 VSUBS 0.047f
C4320 VOUT.t510 VSUBS 0.0294f
C4321 VOUT.t454 VSUBS 0.0294f
C4322 VOUT.n197 VSUBS 0.0711f
C4323 VOUT.n198 VSUBS 0.0264f
C4324 VOUT.n199 VSUBS 0.071f
C4325 VOUT.n200 VSUBS 0.0182f
C4326 VOUT.n201 VSUBS 0.0089f
C4327 VOUT.n202 VSUBS 0.029f
C4328 VOUT.n203 VSUBS 0.22f
C4329 VOUT.n204 VSUBS 0.226f
C4330 VOUT.n205 VSUBS 0.047f
C4331 VOUT.t456 VSUBS 0.0294f
C4332 VOUT.t14 VSUBS 0.0294f
C4333 VOUT.n206 VSUBS 0.0711f
C4334 VOUT.n207 VSUBS 0.0264f
C4335 VOUT.n208 VSUBS 0.071f
C4336 VOUT.n209 VSUBS 0.0182f
C4337 VOUT.n210 VSUBS 0.0089f
C4338 VOUT.n211 VSUBS 0.029f
C4339 VOUT.n212 VSUBS 0.22f
C4340 VOUT.n213 VSUBS 0.226f
C4341 VOUT.n214 VSUBS 0.047f
C4342 VOUT.t396 VSUBS 0.0294f
C4343 VOUT.t97 VSUBS 0.0294f
C4344 VOUT.n215 VSUBS 0.0711f
C4345 VOUT.n216 VSUBS 0.0264f
C4346 VOUT.n217 VSUBS 0.071f
C4347 VOUT.n218 VSUBS 0.0182f
C4348 VOUT.n219 VSUBS 0.0089f
C4349 VOUT.n220 VSUBS 0.029f
C4350 VOUT.n221 VSUBS 0.22f
C4351 VOUT.n222 VSUBS 0.226f
C4352 VOUT.n223 VSUBS 0.047f
C4353 VOUT.t339 VSUBS 0.0294f
C4354 VOUT.t436 VSUBS 0.0294f
C4355 VOUT.n224 VSUBS 0.0711f
C4356 VOUT.n225 VSUBS 0.0264f
C4357 VOUT.n226 VSUBS 0.071f
C4358 VOUT.n227 VSUBS 0.0182f
C4359 VOUT.n228 VSUBS 0.0089f
C4360 VOUT.n229 VSUBS 0.029f
C4361 VOUT.n230 VSUBS 0.22f
C4362 VOUT.n231 VSUBS 0.226f
C4363 VOUT.n232 VSUBS 0.047f
C4364 VOUT.t517 VSUBS 0.0294f
C4365 VOUT.t341 VSUBS 0.0294f
C4366 VOUT.n233 VSUBS 0.0711f
C4367 VOUT.n234 VSUBS 0.0264f
C4368 VOUT.n235 VSUBS 0.071f
C4369 VOUT.n236 VSUBS 0.0182f
C4370 VOUT.n237 VSUBS 0.0089f
C4371 VOUT.n238 VSUBS 0.029f
C4372 VOUT.n239 VSUBS 0.22f
C4373 VOUT.n240 VSUBS 0.226f
C4374 VOUT.n241 VSUBS 0.047f
C4375 VOUT.t417 VSUBS 0.0294f
C4376 VOUT.t445 VSUBS 0.0294f
C4377 VOUT.n242 VSUBS 0.0711f
C4378 VOUT.n243 VSUBS 0.0264f
C4379 VOUT.n244 VSUBS 0.071f
C4380 VOUT.n245 VSUBS 0.0182f
C4381 VOUT.n246 VSUBS 0.0089f
C4382 VOUT.n247 VSUBS 0.029f
C4383 VOUT.n248 VSUBS 0.22f
C4384 VOUT.n249 VSUBS 0.226f
C4385 VOUT.n250 VSUBS 0.047f
C4386 VOUT.t434 VSUBS 0.0294f
C4387 VOUT.t380 VSUBS 0.0294f
C4388 VOUT.n251 VSUBS 0.0711f
C4389 VOUT.n252 VSUBS 0.0264f
C4390 VOUT.n253 VSUBS 0.071f
C4391 VOUT.n254 VSUBS 0.0182f
C4392 VOUT.n255 VSUBS 0.0089f
C4393 VOUT.n256 VSUBS 0.029f
C4394 VOUT.n257 VSUBS 0.22f
C4395 VOUT.n258 VSUBS 0.226f
C4396 VOUT.n259 VSUBS 0.047f
C4397 VOUT.t359 VSUBS 0.0294f
C4398 VOUT.t433 VSUBS 0.0294f
C4399 VOUT.n260 VSUBS 0.0711f
C4400 VOUT.n261 VSUBS 0.0264f
C4401 VOUT.n262 VSUBS 0.071f
C4402 VOUT.n263 VSUBS 0.0182f
C4403 VOUT.n264 VSUBS 0.0089f
C4404 VOUT.n265 VSUBS 0.029f
C4405 VOUT.n266 VSUBS 0.22f
C4406 VOUT.n267 VSUBS 0.226f
C4407 VOUT.n268 VSUBS 0.047f
C4408 VOUT.t457 VSUBS 0.0294f
C4409 VOUT.t420 VSUBS 0.0294f
C4410 VOUT.n269 VSUBS 0.0711f
C4411 VOUT.n270 VSUBS 0.0264f
C4412 VOUT.n271 VSUBS 0.071f
C4413 VOUT.n272 VSUBS 0.0182f
C4414 VOUT.n273 VSUBS 0.0089f
C4415 VOUT.n274 VSUBS 0.029f
C4416 VOUT.n275 VSUBS 0.22f
C4417 VOUT.n276 VSUBS 0.226f
C4418 VOUT.n277 VSUBS 0.047f
C4419 VOUT.t128 VSUBS 0.0294f
C4420 VOUT.t28 VSUBS 0.0294f
C4421 VOUT.n278 VSUBS 0.0711f
C4422 VOUT.n279 VSUBS 0.0264f
C4423 VOUT.n280 VSUBS 0.071f
C4424 VOUT.n281 VSUBS 0.0182f
C4425 VOUT.n282 VSUBS 0.0089f
C4426 VOUT.n283 VSUBS 0.029f
C4427 VOUT.n284 VSUBS 0.22f
C4428 VOUT.n285 VSUBS 0.226f
C4429 VOUT.n286 VSUBS 0.047f
C4430 VOUT.t515 VSUBS 0.0294f
C4431 VOUT.t60 VSUBS 0.0294f
C4432 VOUT.n287 VSUBS 0.0711f
C4433 VOUT.n288 VSUBS 0.0264f
C4434 VOUT.n289 VSUBS 0.071f
C4435 VOUT.n290 VSUBS 0.0182f
C4436 VOUT.n291 VSUBS 0.0089f
C4437 VOUT.n292 VSUBS 0.029f
C4438 VOUT.n293 VSUBS 0.22f
C4439 VOUT.n294 VSUBS 0.226f
C4440 VOUT.n295 VSUBS 0.047f
C4441 VOUT.t36 VSUBS 0.0294f
C4442 VOUT.t432 VSUBS 0.0294f
C4443 VOUT.n296 VSUBS 0.0711f
C4444 VOUT.n297 VSUBS 0.0264f
C4445 VOUT.n298 VSUBS 0.071f
C4446 VOUT.n299 VSUBS 0.0182f
C4447 VOUT.n300 VSUBS 0.0089f
C4448 VOUT.n301 VSUBS 0.029f
C4449 VOUT.n302 VSUBS 0.22f
C4450 VOUT.n303 VSUBS 0.226f
C4451 VOUT.n304 VSUBS 0.047f
C4452 VOUT.t69 VSUBS 0.0294f
C4453 VOUT.t346 VSUBS 0.0294f
C4454 VOUT.n305 VSUBS 0.0711f
C4455 VOUT.n306 VSUBS 0.0264f
C4456 VOUT.n307 VSUBS 0.071f
C4457 VOUT.n308 VSUBS 0.0182f
C4458 VOUT.n309 VSUBS 0.0089f
C4459 VOUT.n310 VSUBS 0.029f
C4460 VOUT.n311 VSUBS 0.22f
C4461 VOUT.n312 VSUBS 0.226f
C4462 VOUT.n313 VSUBS 0.047f
C4463 VOUT.t516 VSUBS 0.0294f
C4464 VOUT.t408 VSUBS 0.0294f
C4465 VOUT.n314 VSUBS 0.0711f
C4466 VOUT.n315 VSUBS 0.0264f
C4467 VOUT.n316 VSUBS 0.071f
C4468 VOUT.n317 VSUBS 0.0182f
C4469 VOUT.n318 VSUBS 0.0089f
C4470 VOUT.n319 VSUBS 0.029f
C4471 VOUT.n320 VSUBS 0.22f
C4472 VOUT.n321 VSUBS 0.226f
C4473 VOUT.n322 VSUBS 0.047f
C4474 VOUT.t33 VSUBS 0.0294f
C4475 VOUT.t54 VSUBS 0.0294f
C4476 VOUT.n323 VSUBS 0.0711f
C4477 VOUT.n324 VSUBS 0.0264f
C4478 VOUT.n325 VSUBS 0.071f
C4479 VOUT.n326 VSUBS 0.0182f
C4480 VOUT.n327 VSUBS 0.0089f
C4481 VOUT.n328 VSUBS 0.029f
C4482 VOUT.n329 VSUBS 0.22f
C4483 VOUT.n330 VSUBS 0.226f
C4484 VOUT.n331 VSUBS 0.047f
C4485 VOUT.t480 VSUBS 0.0294f
C4486 VOUT.t137 VSUBS 0.0294f
C4487 VOUT.n332 VSUBS 0.0711f
C4488 VOUT.n333 VSUBS 0.0264f
C4489 VOUT.n334 VSUBS 0.071f
C4490 VOUT.n335 VSUBS 0.0182f
C4491 VOUT.n336 VSUBS 0.0089f
C4492 VOUT.n337 VSUBS 0.029f
C4493 VOUT.n338 VSUBS 0.22f
C4494 VOUT.n339 VSUBS 0.226f
C4495 VOUT.n340 VSUBS 0.047f
C4496 VOUT.t409 VSUBS 0.0294f
C4497 VOUT.t416 VSUBS 0.0294f
C4498 VOUT.n341 VSUBS 0.0711f
C4499 VOUT.n342 VSUBS 0.0264f
C4500 VOUT.n343 VSUBS 0.071f
C4501 VOUT.n344 VSUBS 0.0182f
C4502 VOUT.n345 VSUBS 0.0089f
C4503 VOUT.n346 VSUBS 0.029f
C4504 VOUT.n347 VSUBS 0.22f
C4505 VOUT.n348 VSUBS 0.226f
C4506 VOUT.n349 VSUBS 0.047f
C4507 VOUT.t443 VSUBS 0.0294f
C4508 VOUT.t135 VSUBS 0.0294f
C4509 VOUT.n350 VSUBS 0.0711f
C4510 VOUT.n351 VSUBS 0.0264f
C4511 VOUT.n352 VSUBS 0.071f
C4512 VOUT.n353 VSUBS 0.0182f
C4513 VOUT.n354 VSUBS 0.0089f
C4514 VOUT.n355 VSUBS 0.029f
C4515 VOUT.n356 VSUBS 0.22f
C4516 VOUT.n357 VSUBS 0.226f
C4517 VOUT.n358 VSUBS 0.047f
C4518 VOUT.t403 VSUBS 0.0294f
C4519 VOUT.t43 VSUBS 0.0294f
C4520 VOUT.n359 VSUBS 0.0711f
C4521 VOUT.n360 VSUBS 0.0264f
C4522 VOUT.n361 VSUBS 0.071f
C4523 VOUT.n362 VSUBS 0.0182f
C4524 VOUT.n363 VSUBS 0.0089f
C4525 VOUT.n364 VSUBS 0.029f
C4526 VOUT.n365 VSUBS 0.22f
C4527 VOUT.n366 VSUBS 0.226f
C4528 VOUT.n367 VSUBS 0.047f
C4529 VOUT.t518 VSUBS 0.0294f
C4530 VOUT.n368 VSUBS 0.1f
C4531 VOUT.n369 VSUBS 0.0264f
C4532 VOUT.n370 VSUBS 0.071f
C4533 VOUT.n371 VSUBS 0.0182f
C4534 VOUT.n372 VSUBS 0.0089f
C4535 VOUT.n373 VSUBS 0.029f
C4536 VOUT.n374 VSUBS 0.22f
C4537 VOUT.n375 VSUBS 0.113f
C4538 VOUT.n376 VSUBS 0.047f
C4539 VOUT.t475 VSUBS 0.0294f
C4540 VOUT.n377 VSUBS 0.1f
C4541 VOUT.n378 VSUBS 0.0264f
C4542 VOUT.n379 VSUBS 0.071f
C4543 VOUT.n380 VSUBS 0.0182f
C4544 VOUT.n381 VSUBS 0.0089f
C4545 VOUT.n382 VSUBS 0.034f
C4546 VOUT.n383 VSUBS 0.322f
C4547 VOUT.n384 VSUBS 0.047f
C4548 VOUT.t470 VSUBS 0.0294f
C4549 VOUT.t461 VSUBS 0.0294f
C4550 VOUT.n385 VSUBS 0.0711f
C4551 VOUT.n386 VSUBS 0.0264f
C4552 VOUT.n387 VSUBS 0.071f
C4553 VOUT.n388 VSUBS 0.0182f
C4554 VOUT.n389 VSUBS 0.0089f
C4555 VOUT.n390 VSUBS 0.029f
C4556 VOUT.n391 VSUBS 0.22f
C4557 VOUT.n392 VSUBS 0.226f
C4558 VOUT.n393 VSUBS 0.047f
C4559 VOUT.t476 VSUBS 0.0294f
C4560 VOUT.t398 VSUBS 0.0294f
C4561 VOUT.n394 VSUBS 0.0711f
C4562 VOUT.n395 VSUBS 0.0264f
C4563 VOUT.n396 VSUBS 0.071f
C4564 VOUT.n397 VSUBS 0.0182f
C4565 VOUT.n398 VSUBS 0.0089f
C4566 VOUT.n399 VSUBS 0.029f
C4567 VOUT.n400 VSUBS 0.22f
C4568 VOUT.n401 VSUBS 0.226f
C4569 VOUT.n402 VSUBS 0.047f
C4570 VOUT.t360 VSUBS 0.0294f
C4571 VOUT.t38 VSUBS 0.0294f
C4572 VOUT.n403 VSUBS 0.0711f
C4573 VOUT.n404 VSUBS 0.0264f
C4574 VOUT.n405 VSUBS 0.071f
C4575 VOUT.n406 VSUBS 0.0182f
C4576 VOUT.n407 VSUBS 0.0089f
C4577 VOUT.n408 VSUBS 0.029f
C4578 VOUT.n409 VSUBS 0.22f
C4579 VOUT.n410 VSUBS 0.226f
C4580 VOUT.n411 VSUBS 0.047f
C4581 VOUT.t467 VSUBS 0.0294f
C4582 VOUT.t11 VSUBS 0.0294f
C4583 VOUT.n412 VSUBS 0.0711f
C4584 VOUT.n413 VSUBS 0.0264f
C4585 VOUT.n414 VSUBS 0.071f
C4586 VOUT.n415 VSUBS 0.0182f
C4587 VOUT.n416 VSUBS 0.0089f
C4588 VOUT.n417 VSUBS 0.029f
C4589 VOUT.n418 VSUBS 0.22f
C4590 VOUT.n419 VSUBS 0.226f
C4591 VOUT.n420 VSUBS 0.047f
C4592 VOUT.t55 VSUBS 0.0294f
C4593 VOUT.t439 VSUBS 0.0294f
C4594 VOUT.n421 VSUBS 0.0711f
C4595 VOUT.n422 VSUBS 0.0264f
C4596 VOUT.n423 VSUBS 0.071f
C4597 VOUT.n424 VSUBS 0.0182f
C4598 VOUT.n425 VSUBS 0.0089f
C4599 VOUT.n426 VSUBS 0.029f
C4600 VOUT.n427 VSUBS 0.22f
C4601 VOUT.n428 VSUBS 0.226f
C4602 VOUT.n429 VSUBS 0.047f
C4603 VOUT.t345 VSUBS 0.0294f
C4604 VOUT.t458 VSUBS 0.0294f
C4605 VOUT.n430 VSUBS 0.0711f
C4606 VOUT.n431 VSUBS 0.0264f
C4607 VOUT.n432 VSUBS 0.071f
C4608 VOUT.n433 VSUBS 0.0182f
C4609 VOUT.n434 VSUBS 0.0089f
C4610 VOUT.n435 VSUBS 0.029f
C4611 VOUT.n436 VSUBS 0.22f
C4612 VOUT.n437 VSUBS 0.226f
C4613 VOUT.n438 VSUBS 0.047f
C4614 VOUT.t450 VSUBS 0.0294f
C4615 VOUT.t15 VSUBS 0.0294f
C4616 VOUT.n439 VSUBS 0.0711f
C4617 VOUT.n440 VSUBS 0.0264f
C4618 VOUT.n441 VSUBS 0.071f
C4619 VOUT.n442 VSUBS 0.0182f
C4620 VOUT.n443 VSUBS 0.0089f
C4621 VOUT.n444 VSUBS 0.029f
C4622 VOUT.n445 VSUBS 0.22f
C4623 VOUT.n446 VSUBS 0.226f
C4624 VOUT.n447 VSUBS 0.047f
C4625 VOUT.t474 VSUBS 0.0294f
C4626 VOUT.t401 VSUBS 0.0294f
C4627 VOUT.n448 VSUBS 0.0711f
C4628 VOUT.n449 VSUBS 0.0264f
C4629 VOUT.n450 VSUBS 0.071f
C4630 VOUT.n451 VSUBS 0.0182f
C4631 VOUT.n452 VSUBS 0.0089f
C4632 VOUT.n453 VSUBS 0.029f
C4633 VOUT.n454 VSUBS 0.22f
C4634 VOUT.n455 VSUBS 0.226f
C4635 VOUT.n456 VSUBS 0.047f
C4636 VOUT.t455 VSUBS 0.0294f
C4637 VOUT.t348 VSUBS 0.0294f
C4638 VOUT.n457 VSUBS 0.0711f
C4639 VOUT.n458 VSUBS 0.0264f
C4640 VOUT.n459 VSUBS 0.071f
C4641 VOUT.n460 VSUBS 0.0182f
C4642 VOUT.n461 VSUBS 0.0089f
C4643 VOUT.n462 VSUBS 0.029f
C4644 VOUT.n463 VSUBS 0.22f
C4645 VOUT.n464 VSUBS 0.226f
C4646 VOUT.n465 VSUBS 0.047f
C4647 VOUT.t442 VSUBS 0.0294f
C4648 VOUT.t6 VSUBS 0.0294f
C4649 VOUT.n466 VSUBS 0.0711f
C4650 VOUT.n467 VSUBS 0.0264f
C4651 VOUT.n468 VSUBS 0.071f
C4652 VOUT.n469 VSUBS 0.0182f
C4653 VOUT.n470 VSUBS 0.0089f
C4654 VOUT.n471 VSUBS 0.029f
C4655 VOUT.n472 VSUBS 0.22f
C4656 VOUT.n473 VSUBS 0.226f
C4657 VOUT.n474 VSUBS 0.047f
C4658 VOUT.t446 VSUBS 0.0294f
C4659 VOUT.t138 VSUBS 0.0294f
C4660 VOUT.n475 VSUBS 0.0711f
C4661 VOUT.n476 VSUBS 0.0264f
C4662 VOUT.n477 VSUBS 0.071f
C4663 VOUT.n478 VSUBS 0.0182f
C4664 VOUT.n479 VSUBS 0.0089f
C4665 VOUT.n480 VSUBS 0.029f
C4666 VOUT.n481 VSUBS 0.22f
C4667 VOUT.n482 VSUBS 0.226f
C4668 VOUT.n483 VSUBS 0.047f
C4669 VOUT.t511 VSUBS 0.0294f
C4670 VOUT.t471 VSUBS 0.0294f
C4671 VOUT.n484 VSUBS 0.0711f
C4672 VOUT.n485 VSUBS 0.0264f
C4673 VOUT.n486 VSUBS 0.071f
C4674 VOUT.n487 VSUBS 0.0182f
C4675 VOUT.n488 VSUBS 0.0089f
C4676 VOUT.n489 VSUBS 0.029f
C4677 VOUT.n490 VSUBS 0.22f
C4678 VOUT.n491 VSUBS 0.226f
C4679 VOUT.n492 VSUBS 0.047f
C4680 VOUT.t392 VSUBS 0.0294f
C4681 VOUT.t437 VSUBS 0.0294f
C4682 VOUT.n493 VSUBS 0.0711f
C4683 VOUT.n494 VSUBS 0.0264f
C4684 VOUT.n495 VSUBS 0.071f
C4685 VOUT.n496 VSUBS 0.0182f
C4686 VOUT.n497 VSUBS 0.0089f
C4687 VOUT.n498 VSUBS 0.029f
C4688 VOUT.n499 VSUBS 0.22f
C4689 VOUT.n500 VSUBS 0.226f
C4690 VOUT.n501 VSUBS 0.047f
C4691 VOUT.t16 VSUBS 0.0294f
C4692 VOUT.t519 VSUBS 0.0294f
C4693 VOUT.n502 VSUBS 0.0711f
C4694 VOUT.n503 VSUBS 0.0264f
C4695 VOUT.n504 VSUBS 0.071f
C4696 VOUT.n505 VSUBS 0.0182f
C4697 VOUT.n506 VSUBS 0.0089f
C4698 VOUT.n507 VSUBS 0.029f
C4699 VOUT.n508 VSUBS 0.22f
C4700 VOUT.n509 VSUBS 0.226f
C4701 VOUT.n510 VSUBS 0.047f
C4702 VOUT.t7 VSUBS 0.0294f
C4703 VOUT.t399 VSUBS 0.0294f
C4704 VOUT.n511 VSUBS 0.0711f
C4705 VOUT.n512 VSUBS 0.0264f
C4706 VOUT.n513 VSUBS 0.071f
C4707 VOUT.n514 VSUBS 0.0182f
C4708 VOUT.n515 VSUBS 0.0089f
C4709 VOUT.n516 VSUBS 0.029f
C4710 VOUT.n517 VSUBS 0.22f
C4711 VOUT.n518 VSUBS 0.226f
C4712 VOUT.n519 VSUBS 0.047f
C4713 VOUT.t469 VSUBS 0.0294f
C4714 VOUT.t482 VSUBS 0.0294f
C4715 VOUT.n520 VSUBS 0.0711f
C4716 VOUT.n521 VSUBS 0.0264f
C4717 VOUT.n522 VSUBS 0.071f
C4718 VOUT.n523 VSUBS 0.0182f
C4719 VOUT.n524 VSUBS 0.0089f
C4720 VOUT.n525 VSUBS 0.029f
C4721 VOUT.n526 VSUBS 0.22f
C4722 VOUT.n527 VSUBS 0.226f
C4723 VOUT.n528 VSUBS 0.047f
C4724 VOUT.t113 VSUBS 0.0294f
C4725 VOUT.t400 VSUBS 0.0294f
C4726 VOUT.n529 VSUBS 0.0711f
C4727 VOUT.n530 VSUBS 0.0264f
C4728 VOUT.n531 VSUBS 0.071f
C4729 VOUT.n532 VSUBS 0.0182f
C4730 VOUT.n533 VSUBS 0.0089f
C4731 VOUT.n534 VSUBS 0.029f
C4732 VOUT.n535 VSUBS 0.22f
C4733 VOUT.n536 VSUBS 0.226f
C4734 VOUT.n537 VSUBS 0.047f
C4735 VOUT.t453 VSUBS 0.0294f
C4736 VOUT.t1 VSUBS 0.0294f
C4737 VOUT.n538 VSUBS 0.0711f
C4738 VOUT.n539 VSUBS 0.0264f
C4739 VOUT.n540 VSUBS 0.071f
C4740 VOUT.n541 VSUBS 0.0182f
C4741 VOUT.n542 VSUBS 0.0089f
C4742 VOUT.n543 VSUBS 0.029f
C4743 VOUT.n544 VSUBS 0.22f
C4744 VOUT.n545 VSUBS 0.226f
C4745 VOUT.n546 VSUBS 0.047f
C4746 VOUT.t468 VSUBS 0.0294f
C4747 VOUT.t411 VSUBS 0.0294f
C4748 VOUT.n547 VSUBS 0.0711f
C4749 VOUT.n548 VSUBS 0.0264f
C4750 VOUT.n549 VSUBS 0.071f
C4751 VOUT.n550 VSUBS 0.0182f
C4752 VOUT.n551 VSUBS 0.0089f
C4753 VOUT.n552 VSUBS 0.029f
C4754 VOUT.n553 VSUBS 0.22f
C4755 VOUT.n554 VSUBS 0.226f
C4756 VOUT.n555 VSUBS 0.047f
C4757 VOUT.t460 VSUBS 0.0294f
C4758 VOUT.n556 VSUBS 0.1f
C4759 VOUT.n557 VSUBS 0.0264f
C4760 VOUT.n558 VSUBS 0.071f
C4761 VOUT.n559 VSUBS 0.0182f
C4762 VOUT.n560 VSUBS 0.0089f
C4763 VOUT.n561 VSUBS 0.029f
C4764 VOUT.n562 VSUBS 0.22f
C4765 VOUT.n563 VSUBS 0.679f
C4766 VOUT.n564 VSUBS 1.41f
C4767 VOUT.n565 VSUBS 1.98f
C4768 VOUT.t253 VSUBS 0.0294f
C4769 VOUT.n566 VSUBS 0.0983f
C4770 VOUT.n567 VSUBS 0.0312f
C4771 VOUT.n568 VSUBS 0.041f
C4772 VOUT.n569 VSUBS 0.0646f
C4773 VOUT.n570 VSUBS 0.0191f
C4774 VOUT.n571 VSUBS 0.00957f
C4775 VOUT.n572 VSUBS 0.0373f
C4776 VOUT.n573 VSUBS 0.322f
C4777 VOUT.n574 VSUBS 0.223f
C4778 VOUT.t153 VSUBS 0.0294f
C4779 VOUT.t306 VSUBS 0.0294f
C4780 VOUT.n575 VSUBS 0.069f
C4781 VOUT.n576 VSUBS 0.0312f
C4782 VOUT.n577 VSUBS 0.0365f
C4783 VOUT.n578 VSUBS 0.0646f
C4784 VOUT.n579 VSUBS 0.0191f
C4785 VOUT.n580 VSUBS 0.00957f
C4786 VOUT.n581 VSUBS 0.0373f
C4787 VOUT.n582 VSUBS 0.223f
C4788 VOUT.n583 VSUBS 0.223f
C4789 VOUT.t286 VSUBS 0.0294f
C4790 VOUT.t235 VSUBS 0.0294f
C4791 VOUT.n584 VSUBS 0.069f
C4792 VOUT.n585 VSUBS 0.0312f
C4793 VOUT.n586 VSUBS 0.0365f
C4794 VOUT.n587 VSUBS 0.0646f
C4795 VOUT.n588 VSUBS 0.0191f
C4796 VOUT.n589 VSUBS 0.00957f
C4797 VOUT.n590 VSUBS 0.0373f
C4798 VOUT.n591 VSUBS 0.223f
C4799 VOUT.n592 VSUBS 0.223f
C4800 VOUT.t180 VSUBS 0.0294f
C4801 VOUT.t334 VSUBS 0.0294f
C4802 VOUT.n593 VSUBS 0.069f
C4803 VOUT.n594 VSUBS 0.0312f
C4804 VOUT.n595 VSUBS 0.0365f
C4805 VOUT.n596 VSUBS 0.0646f
C4806 VOUT.n597 VSUBS 0.0191f
C4807 VOUT.n598 VSUBS 0.00957f
C4808 VOUT.n599 VSUBS 0.0373f
C4809 VOUT.n600 VSUBS 0.223f
C4810 VOUT.n601 VSUBS 0.223f
C4811 VOUT.t183 VSUBS 0.0294f
C4812 VOUT.t284 VSUBS 0.0294f
C4813 VOUT.n602 VSUBS 0.069f
C4814 VOUT.n603 VSUBS 0.0312f
C4815 VOUT.n604 VSUBS 0.0365f
C4816 VOUT.n605 VSUBS 0.0646f
C4817 VOUT.n606 VSUBS 0.0191f
C4818 VOUT.n607 VSUBS 0.00957f
C4819 VOUT.n608 VSUBS 0.0373f
C4820 VOUT.n609 VSUBS 0.223f
C4821 VOUT.n610 VSUBS 0.223f
C4822 VOUT.t263 VSUBS 0.0294f
C4823 VOUT.t216 VSUBS 0.0294f
C4824 VOUT.n611 VSUBS 0.069f
C4825 VOUT.n612 VSUBS 0.0312f
C4826 VOUT.n613 VSUBS 0.0365f
C4827 VOUT.n614 VSUBS 0.0646f
C4828 VOUT.n615 VSUBS 0.0191f
C4829 VOUT.n616 VSUBS 0.00957f
C4830 VOUT.n617 VSUBS 0.0373f
C4831 VOUT.n618 VSUBS 0.223f
C4832 VOUT.n619 VSUBS 0.223f
C4833 VOUT.t161 VSUBS 0.0294f
C4834 VOUT.t316 VSUBS 0.0294f
C4835 VOUT.n620 VSUBS 0.069f
C4836 VOUT.n621 VSUBS 0.0312f
C4837 VOUT.n622 VSUBS 0.0365f
C4838 VOUT.n623 VSUBS 0.0646f
C4839 VOUT.n624 VSUBS 0.0191f
C4840 VOUT.n625 VSUBS 0.00957f
C4841 VOUT.n626 VSUBS 0.0373f
C4842 VOUT.n627 VSUBS 0.223f
C4843 VOUT.n628 VSUBS 0.223f
C4844 VOUT.t168 VSUBS 0.0294f
C4845 VOUT.t322 VSUBS 0.0294f
C4846 VOUT.n629 VSUBS 0.069f
C4847 VOUT.n630 VSUBS 0.0312f
C4848 VOUT.n631 VSUBS 0.0365f
C4849 VOUT.n632 VSUBS 0.0646f
C4850 VOUT.n633 VSUBS 0.0191f
C4851 VOUT.n634 VSUBS 0.00957f
C4852 VOUT.n635 VSUBS 0.0373f
C4853 VOUT.n636 VSUBS 0.223f
C4854 VOUT.n637 VSUBS 0.223f
C4855 VOUT.t243 VSUBS 0.0294f
C4856 VOUT.t251 VSUBS 0.0294f
C4857 VOUT.n638 VSUBS 0.069f
C4858 VOUT.n639 VSUBS 0.0312f
C4859 VOUT.n640 VSUBS 0.0365f
C4860 VOUT.n641 VSUBS 0.0646f
C4861 VOUT.n642 VSUBS 0.0191f
C4862 VOUT.n643 VSUBS 0.00957f
C4863 VOUT.n644 VSUBS 0.0373f
C4864 VOUT.n645 VSUBS 0.223f
C4865 VOUT.n646 VSUBS 0.223f
C4866 VOUT.t192 VSUBS 0.0294f
C4867 VOUT.t292 VSUBS 0.0294f
C4868 VOUT.n647 VSUBS 0.069f
C4869 VOUT.n648 VSUBS 0.0312f
C4870 VOUT.n649 VSUBS 0.0365f
C4871 VOUT.n650 VSUBS 0.0646f
C4872 VOUT.n651 VSUBS 0.0191f
C4873 VOUT.n652 VSUBS 0.00957f
C4874 VOUT.n653 VSUBS 0.0373f
C4875 VOUT.n654 VSUBS 0.223f
C4876 VOUT.n655 VSUBS 0.223f
C4877 VOUT.t145 VSUBS 0.0294f
C4878 VOUT.t237 VSUBS 0.0294f
C4879 VOUT.n656 VSUBS 0.069f
C4880 VOUT.n657 VSUBS 0.0312f
C4881 VOUT.n658 VSUBS 0.0365f
C4882 VOUT.n659 VSUBS 0.0646f
C4883 VOUT.n660 VSUBS 0.0191f
C4884 VOUT.n661 VSUBS 0.00957f
C4885 VOUT.n662 VSUBS 0.0373f
C4886 VOUT.n663 VSUBS 0.223f
C4887 VOUT.n664 VSUBS 0.223f
C4888 VOUT.t221 VSUBS 0.0294f
C4889 VOUT.t338 VSUBS 0.0294f
C4890 VOUT.n665 VSUBS 0.069f
C4891 VOUT.n666 VSUBS 0.0312f
C4892 VOUT.n667 VSUBS 0.0365f
C4893 VOUT.n668 VSUBS 0.0646f
C4894 VOUT.n669 VSUBS 0.0191f
C4895 VOUT.n670 VSUBS 0.00957f
C4896 VOUT.n671 VSUBS 0.0373f
C4897 VOUT.n672 VSUBS 0.223f
C4898 VOUT.n673 VSUBS 0.223f
C4899 VOUT.t321 VSUBS 0.0294f
C4900 VOUT.t271 VSUBS 0.0294f
C4901 VOUT.n674 VSUBS 0.069f
C4902 VOUT.n675 VSUBS 0.0312f
C4903 VOUT.n676 VSUBS 0.0365f
C4904 VOUT.n677 VSUBS 0.0646f
C4905 VOUT.n678 VSUBS 0.0191f
C4906 VOUT.n679 VSUBS 0.00957f
C4907 VOUT.n680 VSUBS 0.0373f
C4908 VOUT.n681 VSUBS 0.223f
C4909 VOUT.n682 VSUBS 0.223f
C4910 VOUT.t193 VSUBS 0.0294f
C4911 VOUT.t240 VSUBS 0.0294f
C4912 VOUT.n683 VSUBS 0.069f
C4913 VOUT.n684 VSUBS 0.0312f
C4914 VOUT.n685 VSUBS 0.0365f
C4915 VOUT.n686 VSUBS 0.0646f
C4916 VOUT.n687 VSUBS 0.0191f
C4917 VOUT.n688 VSUBS 0.00957f
C4918 VOUT.n689 VSUBS 0.0373f
C4919 VOUT.n690 VSUBS 0.223f
C4920 VOUT.n691 VSUBS 0.223f
C4921 VOUT.t244 VSUBS 0.0294f
C4922 VOUT.t293 VSUBS 0.0294f
C4923 VOUT.n692 VSUBS 0.069f
C4924 VOUT.n693 VSUBS 0.0312f
C4925 VOUT.n694 VSUBS 0.0365f
C4926 VOUT.n695 VSUBS 0.0646f
C4927 VOUT.n696 VSUBS 0.0191f
C4928 VOUT.n697 VSUBS 0.00957f
C4929 VOUT.n698 VSUBS 0.0373f
C4930 VOUT.n699 VSUBS 0.223f
C4931 VOUT.n700 VSUBS 0.223f
C4932 VOUT.t317 VSUBS 0.0294f
C4933 VOUT.t204 VSUBS 0.0294f
C4934 VOUT.n701 VSUBS 0.069f
C4935 VOUT.n702 VSUBS 0.0312f
C4936 VOUT.n703 VSUBS 0.0365f
C4937 VOUT.n704 VSUBS 0.0646f
C4938 VOUT.n705 VSUBS 0.0191f
C4939 VOUT.n706 VSUBS 0.00957f
C4940 VOUT.n707 VSUBS 0.0373f
C4941 VOUT.n708 VSUBS 0.223f
C4942 VOUT.n709 VSUBS 0.223f
C4943 VOUT.t222 VSUBS 0.0294f
C4944 VOUT.t323 VSUBS 0.0294f
C4945 VOUT.n710 VSUBS 0.069f
C4946 VOUT.n711 VSUBS 0.0312f
C4947 VOUT.n712 VSUBS 0.0365f
C4948 VOUT.n713 VSUBS 0.0646f
C4949 VOUT.n714 VSUBS 0.0191f
C4950 VOUT.n715 VSUBS 0.00957f
C4951 VOUT.n716 VSUBS 0.0373f
C4952 VOUT.n717 VSUBS 0.223f
C4953 VOUT.n718 VSUBS 0.223f
C4954 VOUT.t287 VSUBS 0.0294f
C4955 VOUT.t188 VSUBS 0.0294f
C4956 VOUT.n719 VSUBS 0.069f
C4957 VOUT.n720 VSUBS 0.0312f
C4958 VOUT.n721 VSUBS 0.0365f
C4959 VOUT.n722 VSUBS 0.0646f
C4960 VOUT.n723 VSUBS 0.0191f
C4961 VOUT.n724 VSUBS 0.00957f
C4962 VOUT.n725 VSUBS 0.0373f
C4963 VOUT.n726 VSUBS 0.223f
C4964 VOUT.n727 VSUBS 0.223f
C4965 VOUT.t247 VSUBS 0.0294f
C4966 VOUT.t238 VSUBS 0.0294f
C4967 VOUT.n728 VSUBS 0.069f
C4968 VOUT.n729 VSUBS 0.0312f
C4969 VOUT.n730 VSUBS 0.0365f
C4970 VOUT.n731 VSUBS 0.0646f
C4971 VOUT.n732 VSUBS 0.0191f
C4972 VOUT.n733 VSUBS 0.00957f
C4973 VOUT.n734 VSUBS 0.0373f
C4974 VOUT.n735 VSUBS 0.223f
C4975 VOUT.n736 VSUBS 0.223f
C4976 VOUT.t239 VSUBS 0.0294f
C4977 VOUT.t163 VSUBS 0.0294f
C4978 VOUT.n737 VSUBS 0.069f
C4979 VOUT.n738 VSUBS 0.0312f
C4980 VOUT.n739 VSUBS 0.0365f
C4981 VOUT.n740 VSUBS 0.0646f
C4982 VOUT.n741 VSUBS 0.0191f
C4983 VOUT.n742 VSUBS 0.00957f
C4984 VOUT.n743 VSUBS 0.0373f
C4985 VOUT.n744 VSUBS 0.223f
C4986 VOUT.n745 VSUBS 0.223f
C4987 VOUT.t156 VSUBS 0.0294f
C4988 VOUT.n746 VSUBS 0.0983f
C4989 VOUT.n747 VSUBS 0.0312f
C4990 VOUT.n748 VSUBS 0.0365f
C4991 VOUT.n749 VSUBS 0.0646f
C4992 VOUT.n750 VSUBS 0.0191f
C4993 VOUT.n751 VSUBS 0.00957f
C4994 VOUT.n752 VSUBS 0.0373f
C4995 VOUT.n753 VSUBS 0.119f
C4996 VOUT.t270 VSUBS 0.0294f
C4997 VOUT.n754 VSUBS 0.0983f
C4998 VOUT.n755 VSUBS 0.031f
C4999 VOUT.n756 VSUBS 0.041f
C5000 VOUT.n757 VSUBS 0.0639f
C5001 VOUT.n758 VSUBS 0.0191f
C5002 VOUT.n759 VSUBS 0.00957f
C5003 VOUT.n760 VSUBS 0.0373f
C5004 VOUT.n761 VSUBS 0.322f
C5005 VOUT.n762 VSUBS 0.223f
C5006 VOUT.t165 VSUBS 0.0294f
C5007 VOUT.t319 VSUBS 0.0294f
C5008 VOUT.n763 VSUBS 0.069f
C5009 VOUT.n764 VSUBS 0.031f
C5010 VOUT.n765 VSUBS 0.0365f
C5011 VOUT.n766 VSUBS 0.0639f
C5012 VOUT.n767 VSUBS 0.0191f
C5013 VOUT.n768 VSUBS 0.00957f
C5014 VOUT.n769 VSUBS 0.0373f
C5015 VOUT.n770 VSUBS 0.223f
C5016 VOUT.n771 VSUBS 0.223f
C5017 VOUT.t303 VSUBS 0.0294f
C5018 VOUT.t248 VSUBS 0.0294f
C5019 VOUT.n772 VSUBS 0.069f
C5020 VOUT.n773 VSUBS 0.031f
C5021 VOUT.n774 VSUBS 0.0365f
C5022 VOUT.n775 VSUBS 0.0639f
C5023 VOUT.n776 VSUBS 0.0191f
C5024 VOUT.n777 VSUBS 0.00957f
C5025 VOUT.n778 VSUBS 0.0373f
C5026 VOUT.n779 VSUBS 0.223f
C5027 VOUT.n780 VSUBS 0.223f
C5028 VOUT.t190 VSUBS 0.0294f
C5029 VOUT.t149 VSUBS 0.0294f
C5030 VOUT.n781 VSUBS 0.069f
C5031 VOUT.n782 VSUBS 0.031f
C5032 VOUT.n783 VSUBS 0.0365f
C5033 VOUT.n784 VSUBS 0.0639f
C5034 VOUT.n785 VSUBS 0.0191f
C5035 VOUT.n786 VSUBS 0.00957f
C5036 VOUT.n787 VSUBS 0.0373f
C5037 VOUT.n788 VSUBS 0.223f
C5038 VOUT.n789 VSUBS 0.223f
C5039 VOUT.t195 VSUBS 0.0294f
C5040 VOUT.t302 VSUBS 0.0294f
C5041 VOUT.n790 VSUBS 0.069f
C5042 VOUT.n791 VSUBS 0.031f
C5043 VOUT.n792 VSUBS 0.0365f
C5044 VOUT.n793 VSUBS 0.0639f
C5045 VOUT.n794 VSUBS 0.0191f
C5046 VOUT.n795 VSUBS 0.00957f
C5047 VOUT.n796 VSUBS 0.0373f
C5048 VOUT.n797 VSUBS 0.223f
C5049 VOUT.n798 VSUBS 0.223f
C5050 VOUT.t281 VSUBS 0.0294f
C5051 VOUT.t230 VSUBS 0.0294f
C5052 VOUT.n799 VSUBS 0.069f
C5053 VOUT.n800 VSUBS 0.031f
C5054 VOUT.n801 VSUBS 0.0365f
C5055 VOUT.n802 VSUBS 0.0639f
C5056 VOUT.n803 VSUBS 0.0191f
C5057 VOUT.n804 VSUBS 0.00957f
C5058 VOUT.n805 VSUBS 0.0373f
C5059 VOUT.n806 VSUBS 0.223f
C5060 VOUT.n807 VSUBS 0.223f
C5061 VOUT.t176 VSUBS 0.0294f
C5062 VOUT.t329 VSUBS 0.0294f
C5063 VOUT.n808 VSUBS 0.069f
C5064 VOUT.n809 VSUBS 0.031f
C5065 VOUT.n810 VSUBS 0.0365f
C5066 VOUT.n811 VSUBS 0.0639f
C5067 VOUT.n812 VSUBS 0.0191f
C5068 VOUT.n813 VSUBS 0.00957f
C5069 VOUT.n814 VSUBS 0.0373f
C5070 VOUT.n815 VSUBS 0.223f
C5071 VOUT.n816 VSUBS 0.223f
C5072 VOUT.t181 VSUBS 0.0294f
C5073 VOUT.t336 VSUBS 0.0294f
C5074 VOUT.n817 VSUBS 0.069f
C5075 VOUT.n818 VSUBS 0.031f
C5076 VOUT.n819 VSUBS 0.0365f
C5077 VOUT.n820 VSUBS 0.0639f
C5078 VOUT.n821 VSUBS 0.0191f
C5079 VOUT.n822 VSUBS 0.00957f
C5080 VOUT.n823 VSUBS 0.0373f
C5081 VOUT.n824 VSUBS 0.223f
C5082 VOUT.n825 VSUBS 0.223f
C5083 VOUT.t257 VSUBS 0.0294f
C5084 VOUT.t267 VSUBS 0.0294f
C5085 VOUT.n826 VSUBS 0.069f
C5086 VOUT.n827 VSUBS 0.031f
C5087 VOUT.n828 VSUBS 0.0365f
C5088 VOUT.n829 VSUBS 0.0639f
C5089 VOUT.n830 VSUBS 0.0191f
C5090 VOUT.n831 VSUBS 0.00957f
C5091 VOUT.n832 VSUBS 0.0373f
C5092 VOUT.n833 VSUBS 0.223f
C5093 VOUT.n834 VSUBS 0.223f
C5094 VOUT.t200 VSUBS 0.0294f
C5095 VOUT.t309 VSUBS 0.0294f
C5096 VOUT.n835 VSUBS 0.069f
C5097 VOUT.n836 VSUBS 0.031f
C5098 VOUT.n837 VSUBS 0.0365f
C5099 VOUT.n838 VSUBS 0.0639f
C5100 VOUT.n839 VSUBS 0.0191f
C5101 VOUT.n840 VSUBS 0.00957f
C5102 VOUT.n841 VSUBS 0.0373f
C5103 VOUT.n842 VSUBS 0.223f
C5104 VOUT.n843 VSUBS 0.223f
C5105 VOUT.t159 VSUBS 0.0294f
C5106 VOUT.t252 VSUBS 0.0294f
C5107 VOUT.n844 VSUBS 0.069f
C5108 VOUT.n845 VSUBS 0.031f
C5109 VOUT.n846 VSUBS 0.0365f
C5110 VOUT.n847 VSUBS 0.0639f
C5111 VOUT.n848 VSUBS 0.0191f
C5112 VOUT.n849 VSUBS 0.00957f
C5113 VOUT.n850 VSUBS 0.0373f
C5114 VOUT.n851 VSUBS 0.223f
C5115 VOUT.n852 VSUBS 0.223f
C5116 VOUT.t234 VSUBS 0.0294f
C5117 VOUT.t155 VSUBS 0.0294f
C5118 VOUT.n853 VSUBS 0.069f
C5119 VOUT.n854 VSUBS 0.031f
C5120 VOUT.n855 VSUBS 0.0365f
C5121 VOUT.n856 VSUBS 0.0639f
C5122 VOUT.n857 VSUBS 0.0191f
C5123 VOUT.n858 VSUBS 0.00957f
C5124 VOUT.n859 VSUBS 0.0373f
C5125 VOUT.n860 VSUBS 0.223f
C5126 VOUT.n861 VSUBS 0.223f
C5127 VOUT.t333 VSUBS 0.0294f
C5128 VOUT.t285 VSUBS 0.0294f
C5129 VOUT.n862 VSUBS 0.069f
C5130 VOUT.n863 VSUBS 0.031f
C5131 VOUT.n864 VSUBS 0.0365f
C5132 VOUT.n865 VSUBS 0.0639f
C5133 VOUT.n866 VSUBS 0.0191f
C5134 VOUT.n867 VSUBS 0.00957f
C5135 VOUT.n868 VSUBS 0.0373f
C5136 VOUT.n869 VSUBS 0.223f
C5137 VOUT.n870 VSUBS 0.223f
C5138 VOUT.t201 VSUBS 0.0294f
C5139 VOUT.t256 VSUBS 0.0294f
C5140 VOUT.n871 VSUBS 0.069f
C5141 VOUT.n872 VSUBS 0.031f
C5142 VOUT.n873 VSUBS 0.0365f
C5143 VOUT.n874 VSUBS 0.0639f
C5144 VOUT.n875 VSUBS 0.0191f
C5145 VOUT.n876 VSUBS 0.00957f
C5146 VOUT.n877 VSUBS 0.0373f
C5147 VOUT.n878 VSUBS 0.223f
C5148 VOUT.n879 VSUBS 0.223f
C5149 VOUT.t259 VSUBS 0.0294f
C5150 VOUT.t311 VSUBS 0.0294f
C5151 VOUT.n880 VSUBS 0.069f
C5152 VOUT.n881 VSUBS 0.031f
C5153 VOUT.n882 VSUBS 0.0365f
C5154 VOUT.n883 VSUBS 0.0639f
C5155 VOUT.n884 VSUBS 0.0191f
C5156 VOUT.n885 VSUBS 0.00957f
C5157 VOUT.n886 VSUBS 0.0373f
C5158 VOUT.n887 VSUBS 0.223f
C5159 VOUT.n888 VSUBS 0.223f
C5160 VOUT.t330 VSUBS 0.0294f
C5161 VOUT.t213 VSUBS 0.0294f
C5162 VOUT.n889 VSUBS 0.069f
C5163 VOUT.n890 VSUBS 0.031f
C5164 VOUT.n891 VSUBS 0.0365f
C5165 VOUT.n892 VSUBS 0.0639f
C5166 VOUT.n893 VSUBS 0.0191f
C5167 VOUT.n894 VSUBS 0.00957f
C5168 VOUT.n895 VSUBS 0.0373f
C5169 VOUT.n896 VSUBS 0.223f
C5170 VOUT.n897 VSUBS 0.223f
C5171 VOUT.t236 VSUBS 0.0294f
C5172 VOUT.t337 VSUBS 0.0294f
C5173 VOUT.n898 VSUBS 0.069f
C5174 VOUT.n899 VSUBS 0.031f
C5175 VOUT.n900 VSUBS 0.0365f
C5176 VOUT.n901 VSUBS 0.0639f
C5177 VOUT.n902 VSUBS 0.0191f
C5178 VOUT.n903 VSUBS 0.00957f
C5179 VOUT.n904 VSUBS 0.0373f
C5180 VOUT.n905 VSUBS 0.223f
C5181 VOUT.n906 VSUBS 0.223f
C5182 VOUT.t308 VSUBS 0.0294f
C5183 VOUT.t198 VSUBS 0.0294f
C5184 VOUT.n907 VSUBS 0.069f
C5185 VOUT.n908 VSUBS 0.031f
C5186 VOUT.n909 VSUBS 0.0365f
C5187 VOUT.n910 VSUBS 0.0639f
C5188 VOUT.n911 VSUBS 0.0191f
C5189 VOUT.n912 VSUBS 0.00957f
C5190 VOUT.n913 VSUBS 0.0373f
C5191 VOUT.n914 VSUBS 0.223f
C5192 VOUT.n915 VSUBS 0.223f
C5193 VOUT.t262 VSUBS 0.0294f
C5194 VOUT.t254 VSUBS 0.0294f
C5195 VOUT.n916 VSUBS 0.069f
C5196 VOUT.n917 VSUBS 0.031f
C5197 VOUT.n918 VSUBS 0.0365f
C5198 VOUT.n919 VSUBS 0.0639f
C5199 VOUT.n920 VSUBS 0.0191f
C5200 VOUT.n921 VSUBS 0.00957f
C5201 VOUT.n922 VSUBS 0.0373f
C5202 VOUT.n923 VSUBS 0.223f
C5203 VOUT.n924 VSUBS 0.223f
C5204 VOUT.t255 VSUBS 0.0294f
C5205 VOUT.t179 VSUBS 0.0294f
C5206 VOUT.n925 VSUBS 0.069f
C5207 VOUT.n926 VSUBS 0.031f
C5208 VOUT.n927 VSUBS 0.0365f
C5209 VOUT.n928 VSUBS 0.0639f
C5210 VOUT.n929 VSUBS 0.0191f
C5211 VOUT.n930 VSUBS 0.00957f
C5212 VOUT.n931 VSUBS 0.0373f
C5213 VOUT.n932 VSUBS 0.223f
C5214 VOUT.n933 VSUBS 0.223f
C5215 VOUT.t170 VSUBS 0.0294f
C5216 VOUT.n934 VSUBS 0.0983f
C5217 VOUT.n935 VSUBS 0.031f
C5218 VOUT.n936 VSUBS 0.0365f
C5219 VOUT.n937 VSUBS 0.0639f
C5220 VOUT.n938 VSUBS 0.0191f
C5221 VOUT.n939 VSUBS 0.00957f
C5222 VOUT.n940 VSUBS 0.0373f
C5223 VOUT.n941 VSUBS 0.119f
C5224 VOUT.t283 VSUBS 0.0294f
C5225 VOUT.n942 VSUBS 0.0983f
C5226 VOUT.n943 VSUBS 0.0306f
C5227 VOUT.n944 VSUBS 0.041f
C5228 VOUT.n945 VSUBS 0.0631f
C5229 VOUT.n946 VSUBS 0.0193f
C5230 VOUT.n947 VSUBS 0.00976f
C5231 VOUT.n948 VSUBS 0.0373f
C5232 VOUT.n949 VSUBS 0.322f
C5233 VOUT.n950 VSUBS 0.223f
C5234 VOUT.t178 VSUBS 0.0294f
C5235 VOUT.t332 VSUBS 0.0294f
C5236 VOUT.n951 VSUBS 0.0689f
C5237 VOUT.n952 VSUBS 0.0306f
C5238 VOUT.n953 VSUBS 0.0365f
C5239 VOUT.n954 VSUBS 0.0631f
C5240 VOUT.n955 VSUBS 0.0193f
C5241 VOUT.n956 VSUBS 0.00976f
C5242 VOUT.n957 VSUBS 0.0373f
C5243 VOUT.n958 VSUBS 0.223f
C5244 VOUT.n959 VSUBS 0.223f
C5245 VOUT.t315 VSUBS 0.0294f
C5246 VOUT.t261 VSUBS 0.0294f
C5247 VOUT.n960 VSUBS 0.0689f
C5248 VOUT.n961 VSUBS 0.0306f
C5249 VOUT.n962 VSUBS 0.0365f
C5250 VOUT.n963 VSUBS 0.0631f
C5251 VOUT.n964 VSUBS 0.0193f
C5252 VOUT.n965 VSUBS 0.00976f
C5253 VOUT.n966 VSUBS 0.0373f
C5254 VOUT.n967 VSUBS 0.223f
C5255 VOUT.n968 VSUBS 0.223f
C5256 VOUT.t197 VSUBS 0.0294f
C5257 VOUT.t160 VSUBS 0.0294f
C5258 VOUT.n969 VSUBS 0.0689f
C5259 VOUT.n970 VSUBS 0.0306f
C5260 VOUT.n971 VSUBS 0.0365f
C5261 VOUT.n972 VSUBS 0.0631f
C5262 VOUT.n973 VSUBS 0.0193f
C5263 VOUT.n974 VSUBS 0.00976f
C5264 VOUT.n975 VSUBS 0.0373f
C5265 VOUT.n976 VSUBS 0.223f
C5266 VOUT.n977 VSUBS 0.223f
C5267 VOUT.t203 VSUBS 0.0294f
C5268 VOUT.t314 VSUBS 0.0294f
C5269 VOUT.n978 VSUBS 0.0689f
C5270 VOUT.n979 VSUBS 0.0306f
C5271 VOUT.n980 VSUBS 0.0365f
C5272 VOUT.n981 VSUBS 0.0631f
C5273 VOUT.n982 VSUBS 0.0193f
C5274 VOUT.n983 VSUBS 0.00976f
C5275 VOUT.n984 VSUBS 0.0373f
C5276 VOUT.n985 VSUBS 0.223f
C5277 VOUT.n986 VSUBS 0.223f
C5278 VOUT.t291 VSUBS 0.0294f
C5279 VOUT.t242 VSUBS 0.0294f
C5280 VOUT.n987 VSUBS 0.0689f
C5281 VOUT.n988 VSUBS 0.0306f
C5282 VOUT.n989 VSUBS 0.0365f
C5283 VOUT.n990 VSUBS 0.0631f
C5284 VOUT.n991 VSUBS 0.0193f
C5285 VOUT.n992 VSUBS 0.00976f
C5286 VOUT.n993 VSUBS 0.0373f
C5287 VOUT.n994 VSUBS 0.223f
C5288 VOUT.n995 VSUBS 0.223f
C5289 VOUT.t185 VSUBS 0.0294f
C5290 VOUT.t142 VSUBS 0.0294f
C5291 VOUT.n996 VSUBS 0.0689f
C5292 VOUT.n997 VSUBS 0.0306f
C5293 VOUT.n998 VSUBS 0.0365f
C5294 VOUT.n999 VSUBS 0.0631f
C5295 VOUT.n1000 VSUBS 0.0193f
C5296 VOUT.n1001 VSUBS 0.00976f
C5297 VOUT.n1002 VSUBS 0.0373f
C5298 VOUT.n1003 VSUBS 0.223f
C5299 VOUT.n1004 VSUBS 0.223f
C5300 VOUT.t191 VSUBS 0.0294f
C5301 VOUT.t150 VSUBS 0.0294f
C5302 VOUT.n1005 VSUBS 0.0689f
C5303 VOUT.n1006 VSUBS 0.0306f
C5304 VOUT.n1007 VSUBS 0.0365f
C5305 VOUT.n1008 VSUBS 0.0631f
C5306 VOUT.n1009 VSUBS 0.0193f
C5307 VOUT.n1010 VSUBS 0.00976f
C5308 VOUT.n1011 VSUBS 0.0373f
C5309 VOUT.n1012 VSUBS 0.223f
C5310 VOUT.n1013 VSUBS 0.223f
C5311 VOUT.t275 VSUBS 0.0294f
C5312 VOUT.t282 VSUBS 0.0294f
C5313 VOUT.n1014 VSUBS 0.0689f
C5314 VOUT.n1015 VSUBS 0.0306f
C5315 VOUT.n1016 VSUBS 0.0365f
C5316 VOUT.n1017 VSUBS 0.0631f
C5317 VOUT.n1018 VSUBS 0.0193f
C5318 VOUT.n1019 VSUBS 0.00976f
C5319 VOUT.n1020 VSUBS 0.0373f
C5320 VOUT.n1021 VSUBS 0.223f
C5321 VOUT.n1022 VSUBS 0.223f
C5322 VOUT.t211 VSUBS 0.0294f
C5323 VOUT.t326 VSUBS 0.0294f
C5324 VOUT.n1023 VSUBS 0.0689f
C5325 VOUT.n1024 VSUBS 0.0306f
C5326 VOUT.n1025 VSUBS 0.0365f
C5327 VOUT.n1026 VSUBS 0.0631f
C5328 VOUT.n1027 VSUBS 0.0193f
C5329 VOUT.n1028 VSUBS 0.00976f
C5330 VOUT.n1029 VSUBS 0.0373f
C5331 VOUT.n1030 VSUBS 0.223f
C5332 VOUT.n1031 VSUBS 0.223f
C5333 VOUT.t171 VSUBS 0.0294f
C5334 VOUT.t265 VSUBS 0.0294f
C5335 VOUT.n1032 VSUBS 0.0689f
C5336 VOUT.n1033 VSUBS 0.0306f
C5337 VOUT.n1034 VSUBS 0.0365f
C5338 VOUT.n1035 VSUBS 0.0631f
C5339 VOUT.n1036 VSUBS 0.0193f
C5340 VOUT.n1037 VSUBS 0.00976f
C5341 VOUT.n1038 VSUBS 0.0373f
C5342 VOUT.n1039 VSUBS 0.223f
C5343 VOUT.n1040 VSUBS 0.223f
C5344 VOUT.t246 VSUBS 0.0294f
C5345 VOUT.t162 VSUBS 0.0294f
C5346 VOUT.n1041 VSUBS 0.0689f
C5347 VOUT.n1042 VSUBS 0.0306f
C5348 VOUT.n1043 VSUBS 0.0365f
C5349 VOUT.n1044 VSUBS 0.0631f
C5350 VOUT.n1045 VSUBS 0.0193f
C5351 VOUT.n1046 VSUBS 0.00976f
C5352 VOUT.n1047 VSUBS 0.0373f
C5353 VOUT.n1048 VSUBS 0.223f
C5354 VOUT.n1049 VSUBS 0.223f
C5355 VOUT.t147 VSUBS 0.0294f
C5356 VOUT.t298 VSUBS 0.0294f
C5357 VOUT.n1050 VSUBS 0.0689f
C5358 VOUT.n1051 VSUBS 0.0306f
C5359 VOUT.n1052 VSUBS 0.0365f
C5360 VOUT.n1053 VSUBS 0.0631f
C5361 VOUT.n1054 VSUBS 0.0193f
C5362 VOUT.n1055 VSUBS 0.00976f
C5363 VOUT.n1056 VSUBS 0.0373f
C5364 VOUT.n1057 VSUBS 0.223f
C5365 VOUT.n1058 VSUBS 0.223f
C5366 VOUT.t212 VSUBS 0.0294f
C5367 VOUT.t269 VSUBS 0.0294f
C5368 VOUT.n1059 VSUBS 0.0689f
C5369 VOUT.n1060 VSUBS 0.0306f
C5370 VOUT.n1061 VSUBS 0.0365f
C5371 VOUT.n1062 VSUBS 0.0631f
C5372 VOUT.n1063 VSUBS 0.0193f
C5373 VOUT.n1064 VSUBS 0.00976f
C5374 VOUT.n1065 VSUBS 0.0373f
C5375 VOUT.n1066 VSUBS 0.223f
C5376 VOUT.n1067 VSUBS 0.223f
C5377 VOUT.t276 VSUBS 0.0294f
C5378 VOUT.t327 VSUBS 0.0294f
C5379 VOUT.n1068 VSUBS 0.0689f
C5380 VOUT.n1069 VSUBS 0.0306f
C5381 VOUT.n1070 VSUBS 0.0365f
C5382 VOUT.n1071 VSUBS 0.0631f
C5383 VOUT.n1072 VSUBS 0.0193f
C5384 VOUT.n1073 VSUBS 0.00976f
C5385 VOUT.n1074 VSUBS 0.0373f
C5386 VOUT.n1075 VSUBS 0.223f
C5387 VOUT.n1076 VSUBS 0.223f
C5388 VOUT.t143 VSUBS 0.0294f
C5389 VOUT.t226 VSUBS 0.0294f
C5390 VOUT.n1077 VSUBS 0.0689f
C5391 VOUT.n1078 VSUBS 0.0306f
C5392 VOUT.n1079 VSUBS 0.0365f
C5393 VOUT.n1080 VSUBS 0.0631f
C5394 VOUT.n1081 VSUBS 0.0193f
C5395 VOUT.n1082 VSUBS 0.00976f
C5396 VOUT.n1083 VSUBS 0.0373f
C5397 VOUT.n1084 VSUBS 0.223f
C5398 VOUT.n1085 VSUBS 0.223f
C5399 VOUT.t249 VSUBS 0.0294f
C5400 VOUT.t151 VSUBS 0.0294f
C5401 VOUT.n1086 VSUBS 0.0689f
C5402 VOUT.n1087 VSUBS 0.0306f
C5403 VOUT.n1088 VSUBS 0.0365f
C5404 VOUT.n1089 VSUBS 0.0631f
C5405 VOUT.n1090 VSUBS 0.0193f
C5406 VOUT.n1091 VSUBS 0.00976f
C5407 VOUT.n1092 VSUBS 0.0373f
C5408 VOUT.n1093 VSUBS 0.223f
C5409 VOUT.n1094 VSUBS 0.223f
C5410 VOUT.t320 VSUBS 0.0294f
C5411 VOUT.t209 VSUBS 0.0294f
C5412 VOUT.n1095 VSUBS 0.0689f
C5413 VOUT.n1096 VSUBS 0.0306f
C5414 VOUT.n1097 VSUBS 0.0365f
C5415 VOUT.n1098 VSUBS 0.0631f
C5416 VOUT.n1099 VSUBS 0.0193f
C5417 VOUT.n1100 VSUBS 0.00976f
C5418 VOUT.n1101 VSUBS 0.0373f
C5419 VOUT.n1102 VSUBS 0.223f
C5420 VOUT.n1103 VSUBS 0.223f
C5421 VOUT.t278 VSUBS 0.0294f
C5422 VOUT.t266 VSUBS 0.0294f
C5423 VOUT.n1104 VSUBS 0.0689f
C5424 VOUT.n1105 VSUBS 0.0306f
C5425 VOUT.n1106 VSUBS 0.0365f
C5426 VOUT.n1107 VSUBS 0.0631f
C5427 VOUT.n1108 VSUBS 0.0193f
C5428 VOUT.n1109 VSUBS 0.00976f
C5429 VOUT.n1110 VSUBS 0.0373f
C5430 VOUT.n1111 VSUBS 0.223f
C5431 VOUT.n1112 VSUBS 0.223f
C5432 VOUT.t268 VSUBS 0.0294f
C5433 VOUT.t187 VSUBS 0.0294f
C5434 VOUT.n1113 VSUBS 0.0689f
C5435 VOUT.n1114 VSUBS 0.0306f
C5436 VOUT.n1115 VSUBS 0.0365f
C5437 VOUT.n1116 VSUBS 0.0631f
C5438 VOUT.n1117 VSUBS 0.0193f
C5439 VOUT.n1118 VSUBS 0.00976f
C5440 VOUT.n1119 VSUBS 0.0373f
C5441 VOUT.n1120 VSUBS 0.223f
C5442 VOUT.n1121 VSUBS 0.223f
C5443 VOUT.t182 VSUBS 0.0294f
C5444 VOUT.n1122 VSUBS 0.0983f
C5445 VOUT.n1123 VSUBS 0.0306f
C5446 VOUT.n1124 VSUBS 0.0365f
C5447 VOUT.n1125 VSUBS 0.0631f
C5448 VOUT.n1126 VSUBS 0.0193f
C5449 VOUT.n1127 VSUBS 0.00976f
C5450 VOUT.n1128 VSUBS 0.0373f
C5451 VOUT.n1129 VSUBS 0.119f
C5452 VOUT.t231 VSUBS 0.0294f
C5453 VOUT.n1130 VSUBS 0.0983f
C5454 VOUT.n1131 VSUBS 0.0304f
C5455 VOUT.n1132 VSUBS 0.041f
C5456 VOUT.n1133 VSUBS 0.0623f
C5457 VOUT.n1134 VSUBS 0.0193f
C5458 VOUT.n1135 VSUBS 0.00976f
C5459 VOUT.n1136 VSUBS 0.0373f
C5460 VOUT.n1137 VSUBS 0.322f
C5461 VOUT.n1138 VSUBS 0.223f
C5462 VOUT.t331 VSUBS 0.0294f
C5463 VOUT.t280 VSUBS 0.0294f
C5464 VOUT.n1139 VSUBS 0.0689f
C5465 VOUT.n1140 VSUBS 0.0304f
C5466 VOUT.n1141 VSUBS 0.0365f
C5467 VOUT.n1142 VSUBS 0.0623f
C5468 VOUT.n1143 VSUBS 0.0193f
C5469 VOUT.n1144 VSUBS 0.00976f
C5470 VOUT.n1145 VSUBS 0.0373f
C5471 VOUT.n1146 VSUBS 0.223f
C5472 VOUT.n1147 VSUBS 0.223f
C5473 VOUT.t260 VSUBS 0.0294f
C5474 VOUT.t214 VSUBS 0.0294f
C5475 VOUT.n1148 VSUBS 0.0689f
C5476 VOUT.n1149 VSUBS 0.0304f
C5477 VOUT.n1150 VSUBS 0.0365f
C5478 VOUT.n1151 VSUBS 0.0623f
C5479 VOUT.n1152 VSUBS 0.0193f
C5480 VOUT.n1153 VSUBS 0.00976f
C5481 VOUT.n1154 VSUBS 0.0373f
C5482 VOUT.n1155 VSUBS 0.223f
C5483 VOUT.n1156 VSUBS 0.223f
C5484 VOUT.t157 VSUBS 0.0294f
C5485 VOUT.t312 VSUBS 0.0294f
C5486 VOUT.n1157 VSUBS 0.0689f
C5487 VOUT.n1158 VSUBS 0.0304f
C5488 VOUT.n1159 VSUBS 0.0365f
C5489 VOUT.n1160 VSUBS 0.0623f
C5490 VOUT.n1161 VSUBS 0.0193f
C5491 VOUT.n1162 VSUBS 0.00976f
C5492 VOUT.n1163 VSUBS 0.0373f
C5493 VOUT.n1164 VSUBS 0.223f
C5494 VOUT.n1165 VSUBS 0.223f
C5495 VOUT.t164 VSUBS 0.0294f
C5496 VOUT.t258 VSUBS 0.0294f
C5497 VOUT.n1166 VSUBS 0.0689f
C5498 VOUT.n1167 VSUBS 0.0304f
C5499 VOUT.n1168 VSUBS 0.0365f
C5500 VOUT.n1169 VSUBS 0.0623f
C5501 VOUT.n1170 VSUBS 0.0193f
C5502 VOUT.n1171 VSUBS 0.00976f
C5503 VOUT.n1172 VSUBS 0.0373f
C5504 VOUT.n1173 VSUBS 0.223f
C5505 VOUT.n1174 VSUBS 0.223f
C5506 VOUT.t241 VSUBS 0.0294f
C5507 VOUT.t202 VSUBS 0.0294f
C5508 VOUT.n1175 VSUBS 0.0689f
C5509 VOUT.n1176 VSUBS 0.0304f
C5510 VOUT.n1177 VSUBS 0.0365f
C5511 VOUT.n1178 VSUBS 0.0623f
C5512 VOUT.n1179 VSUBS 0.0193f
C5513 VOUT.n1180 VSUBS 0.00976f
C5514 VOUT.n1181 VSUBS 0.0373f
C5515 VOUT.n1182 VSUBS 0.223f
C5516 VOUT.n1183 VSUBS 0.223f
C5517 VOUT.t139 VSUBS 0.0294f
C5518 VOUT.t288 VSUBS 0.0294f
C5519 VOUT.n1184 VSUBS 0.0689f
C5520 VOUT.n1185 VSUBS 0.0304f
C5521 VOUT.n1186 VSUBS 0.0365f
C5522 VOUT.n1187 VSUBS 0.0623f
C5523 VOUT.n1188 VSUBS 0.0193f
C5524 VOUT.n1189 VSUBS 0.00976f
C5525 VOUT.n1190 VSUBS 0.0373f
C5526 VOUT.n1191 VSUBS 0.223f
C5527 VOUT.n1192 VSUBS 0.223f
C5528 VOUT.t148 VSUBS 0.0294f
C5529 VOUT.t300 VSUBS 0.0294f
C5530 VOUT.n1193 VSUBS 0.0689f
C5531 VOUT.n1194 VSUBS 0.0304f
C5532 VOUT.n1195 VSUBS 0.0365f
C5533 VOUT.n1196 VSUBS 0.0623f
C5534 VOUT.n1197 VSUBS 0.0193f
C5535 VOUT.n1198 VSUBS 0.00976f
C5536 VOUT.n1199 VSUBS 0.0373f
C5537 VOUT.n1200 VSUBS 0.223f
C5538 VOUT.n1201 VSUBS 0.223f
C5539 VOUT.t223 VSUBS 0.0294f
C5540 VOUT.t229 VSUBS 0.0294f
C5541 VOUT.n1202 VSUBS 0.0689f
C5542 VOUT.n1203 VSUBS 0.0304f
C5543 VOUT.n1204 VSUBS 0.0365f
C5544 VOUT.n1205 VSUBS 0.0623f
C5545 VOUT.n1206 VSUBS 0.0193f
C5546 VOUT.n1207 VSUBS 0.00976f
C5547 VOUT.n1208 VSUBS 0.0373f
C5548 VOUT.n1209 VSUBS 0.223f
C5549 VOUT.n1210 VSUBS 0.223f
C5550 VOUT.t173 VSUBS 0.0294f
C5551 VOUT.t272 VSUBS 0.0294f
C5552 VOUT.n1211 VSUBS 0.0689f
C5553 VOUT.n1212 VSUBS 0.0304f
C5554 VOUT.n1213 VSUBS 0.0365f
C5555 VOUT.n1214 VSUBS 0.0623f
C5556 VOUT.n1215 VSUBS 0.0193f
C5557 VOUT.n1216 VSUBS 0.00976f
C5558 VOUT.n1217 VSUBS 0.0373f
C5559 VOUT.n1218 VSUBS 0.223f
C5560 VOUT.n1219 VSUBS 0.223f
C5561 VOUT.t325 VSUBS 0.0294f
C5562 VOUT.t217 VSUBS 0.0294f
C5563 VOUT.n1220 VSUBS 0.0689f
C5564 VOUT.n1221 VSUBS 0.0304f
C5565 VOUT.n1222 VSUBS 0.0365f
C5566 VOUT.n1223 VSUBS 0.0623f
C5567 VOUT.n1224 VSUBS 0.0193f
C5568 VOUT.n1225 VSUBS 0.00976f
C5569 VOUT.n1226 VSUBS 0.0373f
C5570 VOUT.n1227 VSUBS 0.223f
C5571 VOUT.n1228 VSUBS 0.223f
C5572 VOUT.t206 VSUBS 0.0294f
C5573 VOUT.t318 VSUBS 0.0294f
C5574 VOUT.n1229 VSUBS 0.0689f
C5575 VOUT.n1230 VSUBS 0.0304f
C5576 VOUT.n1231 VSUBS 0.0365f
C5577 VOUT.n1232 VSUBS 0.0623f
C5578 VOUT.n1233 VSUBS 0.0193f
C5579 VOUT.n1234 VSUBS 0.00976f
C5580 VOUT.n1235 VSUBS 0.0373f
C5581 VOUT.n1236 VSUBS 0.223f
C5582 VOUT.n1237 VSUBS 0.223f
C5583 VOUT.t294 VSUBS 0.0294f
C5584 VOUT.t245 VSUBS 0.0294f
C5585 VOUT.n1238 VSUBS 0.0689f
C5586 VOUT.n1239 VSUBS 0.0304f
C5587 VOUT.n1240 VSUBS 0.0365f
C5588 VOUT.n1241 VSUBS 0.0623f
C5589 VOUT.n1242 VSUBS 0.0193f
C5590 VOUT.n1243 VSUBS 0.00976f
C5591 VOUT.n1244 VSUBS 0.0373f
C5592 VOUT.n1245 VSUBS 0.223f
C5593 VOUT.n1246 VSUBS 0.223f
C5594 VOUT.t175 VSUBS 0.0294f
C5595 VOUT.t220 VSUBS 0.0294f
C5596 VOUT.n1247 VSUBS 0.0689f
C5597 VOUT.n1248 VSUBS 0.0304f
C5598 VOUT.n1249 VSUBS 0.0365f
C5599 VOUT.n1250 VSUBS 0.0623f
C5600 VOUT.n1251 VSUBS 0.0193f
C5601 VOUT.n1252 VSUBS 0.00976f
C5602 VOUT.n1253 VSUBS 0.0373f
C5603 VOUT.n1254 VSUBS 0.223f
C5604 VOUT.n1255 VSUBS 0.223f
C5605 VOUT.t224 VSUBS 0.0294f
C5606 VOUT.t273 VSUBS 0.0294f
C5607 VOUT.n1256 VSUBS 0.0689f
C5608 VOUT.n1257 VSUBS 0.0304f
C5609 VOUT.n1258 VSUBS 0.0365f
C5610 VOUT.n1259 VSUBS 0.0623f
C5611 VOUT.n1260 VSUBS 0.0193f
C5612 VOUT.n1261 VSUBS 0.00976f
C5613 VOUT.n1262 VSUBS 0.0373f
C5614 VOUT.n1263 VSUBS 0.223f
C5615 VOUT.n1264 VSUBS 0.223f
C5616 VOUT.t289 VSUBS 0.0294f
C5617 VOUT.t189 VSUBS 0.0294f
C5618 VOUT.n1265 VSUBS 0.0689f
C5619 VOUT.n1266 VSUBS 0.0304f
C5620 VOUT.n1267 VSUBS 0.0365f
C5621 VOUT.n1268 VSUBS 0.0623f
C5622 VOUT.n1269 VSUBS 0.0193f
C5623 VOUT.n1270 VSUBS 0.00976f
C5624 VOUT.n1271 VSUBS 0.0373f
C5625 VOUT.n1272 VSUBS 0.223f
C5626 VOUT.n1273 VSUBS 0.223f
C5627 VOUT.t207 VSUBS 0.0294f
C5628 VOUT.t301 VSUBS 0.0294f
C5629 VOUT.n1274 VSUBS 0.0689f
C5630 VOUT.n1275 VSUBS 0.0304f
C5631 VOUT.n1276 VSUBS 0.0365f
C5632 VOUT.n1277 VSUBS 0.0623f
C5633 VOUT.n1278 VSUBS 0.0193f
C5634 VOUT.n1279 VSUBS 0.00976f
C5635 VOUT.n1280 VSUBS 0.0373f
C5636 VOUT.n1281 VSUBS 0.223f
C5637 VOUT.n1282 VSUBS 0.223f
C5638 VOUT.t264 VSUBS 0.0294f
C5639 VOUT.t169 VSUBS 0.0294f
C5640 VOUT.n1283 VSUBS 0.0689f
C5641 VOUT.n1284 VSUBS 0.0304f
C5642 VOUT.n1285 VSUBS 0.0365f
C5643 VOUT.n1286 VSUBS 0.0623f
C5644 VOUT.n1287 VSUBS 0.0193f
C5645 VOUT.n1288 VSUBS 0.00976f
C5646 VOUT.n1289 VSUBS 0.0373f
C5647 VOUT.n1290 VSUBS 0.223f
C5648 VOUT.n1291 VSUBS 0.223f
C5649 VOUT.t227 VSUBS 0.0294f
C5650 VOUT.t218 VSUBS 0.0294f
C5651 VOUT.n1292 VSUBS 0.0689f
C5652 VOUT.n1293 VSUBS 0.0304f
C5653 VOUT.n1294 VSUBS 0.0365f
C5654 VOUT.n1295 VSUBS 0.0623f
C5655 VOUT.n1296 VSUBS 0.0193f
C5656 VOUT.n1297 VSUBS 0.00976f
C5657 VOUT.n1298 VSUBS 0.0373f
C5658 VOUT.n1299 VSUBS 0.223f
C5659 VOUT.n1300 VSUBS 0.223f
C5660 VOUT.t219 VSUBS 0.0294f
C5661 VOUT.t144 VSUBS 0.0294f
C5662 VOUT.n1301 VSUBS 0.0689f
C5663 VOUT.n1302 VSUBS 0.0304f
C5664 VOUT.n1303 VSUBS 0.0365f
C5665 VOUT.n1304 VSUBS 0.0623f
C5666 VOUT.n1305 VSUBS 0.0193f
C5667 VOUT.n1306 VSUBS 0.00976f
C5668 VOUT.n1307 VSUBS 0.0373f
C5669 VOUT.n1308 VSUBS 0.223f
C5670 VOUT.n1309 VSUBS 0.223f
C5671 VOUT.t335 VSUBS 0.0294f
C5672 VOUT.n1310 VSUBS 0.0983f
C5673 VOUT.n1311 VSUBS 0.0304f
C5674 VOUT.n1312 VSUBS 0.0365f
C5675 VOUT.n1313 VSUBS 0.0623f
C5676 VOUT.n1314 VSUBS 0.0193f
C5677 VOUT.n1315 VSUBS 0.00976f
C5678 VOUT.n1316 VSUBS 0.0373f
C5679 VOUT.n1317 VSUBS 0.119f
C5680 VOUT.t313 VSUBS 0.0294f
C5681 VOUT.n1318 VSUBS 0.0982f
C5682 VOUT.n1319 VSUBS 0.03f
C5683 VOUT.n1320 VSUBS 0.041f
C5684 VOUT.n1321 VSUBS 0.0615f
C5685 VOUT.n1322 VSUBS 0.0195f
C5686 VOUT.n1323 VSUBS 0.00998f
C5687 VOUT.n1324 VSUBS 0.0373f
C5688 VOUT.n1325 VSUBS 0.322f
C5689 VOUT.n1326 VSUBS 0.223f
C5690 VOUT.t196 VSUBS 0.0294f
C5691 VOUT.t158 VSUBS 0.0294f
C5692 VOUT.n1327 VSUBS 0.0689f
C5693 VOUT.n1328 VSUBS 0.03f
C5694 VOUT.n1329 VSUBS 0.0365f
C5695 VOUT.n1330 VSUBS 0.0615f
C5696 VOUT.n1331 VSUBS 0.0195f
C5697 VOUT.n1332 VSUBS 0.00998f
C5698 VOUT.n1333 VSUBS 0.0373f
C5699 VOUT.n1334 VSUBS 0.223f
C5700 VOUT.n1335 VSUBS 0.223f
C5701 VOUT.t141 VSUBS 0.0294f
C5702 VOUT.t290 VSUBS 0.0294f
C5703 VOUT.n1336 VSUBS 0.0689f
C5704 VOUT.n1337 VSUBS 0.03f
C5705 VOUT.n1338 VSUBS 0.0365f
C5706 VOUT.n1339 VSUBS 0.0615f
C5707 VOUT.n1340 VSUBS 0.0195f
C5708 VOUT.n1341 VSUBS 0.00998f
C5709 VOUT.n1342 VSUBS 0.0373f
C5710 VOUT.n1343 VSUBS 0.223f
C5711 VOUT.n1344 VSUBS 0.223f
C5712 VOUT.t215 VSUBS 0.0294f
C5713 VOUT.t184 VSUBS 0.0294f
C5714 VOUT.n1345 VSUBS 0.0689f
C5715 VOUT.n1346 VSUBS 0.03f
C5716 VOUT.n1347 VSUBS 0.0365f
C5717 VOUT.n1348 VSUBS 0.0615f
C5718 VOUT.n1349 VSUBS 0.0195f
C5719 VOUT.n1350 VSUBS 0.00998f
C5720 VOUT.n1351 VSUBS 0.0373f
C5721 VOUT.n1352 VSUBS 0.223f
C5722 VOUT.n1353 VSUBS 0.223f
C5723 VOUT.t225 VSUBS 0.0294f
C5724 VOUT.t140 VSUBS 0.0294f
C5725 VOUT.n1354 VSUBS 0.0689f
C5726 VOUT.n1355 VSUBS 0.03f
C5727 VOUT.n1356 VSUBS 0.0365f
C5728 VOUT.n1357 VSUBS 0.0615f
C5729 VOUT.n1358 VSUBS 0.0195f
C5730 VOUT.n1359 VSUBS 0.00998f
C5731 VOUT.n1360 VSUBS 0.0373f
C5732 VOUT.n1361 VSUBS 0.223f
C5733 VOUT.n1362 VSUBS 0.223f
C5734 VOUT.t324 VSUBS 0.0294f
C5735 VOUT.t274 VSUBS 0.0294f
C5736 VOUT.n1363 VSUBS 0.0689f
C5737 VOUT.n1364 VSUBS 0.03f
C5738 VOUT.n1365 VSUBS 0.0365f
C5739 VOUT.n1366 VSUBS 0.0615f
C5740 VOUT.n1367 VSUBS 0.0195f
C5741 VOUT.n1368 VSUBS 0.00998f
C5742 VOUT.n1369 VSUBS 0.0373f
C5743 VOUT.n1370 VSUBS 0.223f
C5744 VOUT.n1371 VSUBS 0.223f
C5745 VOUT.t205 VSUBS 0.0294f
C5746 VOUT.t166 VSUBS 0.0294f
C5747 VOUT.n1372 VSUBS 0.0689f
C5748 VOUT.n1373 VSUBS 0.03f
C5749 VOUT.n1374 VSUBS 0.0365f
C5750 VOUT.n1375 VSUBS 0.0615f
C5751 VOUT.n1376 VSUBS 0.0195f
C5752 VOUT.n1377 VSUBS 0.00998f
C5753 VOUT.n1378 VSUBS 0.0373f
C5754 VOUT.n1379 VSUBS 0.223f
C5755 VOUT.n1380 VSUBS 0.223f
C5756 VOUT.t210 VSUBS 0.0294f
C5757 VOUT.t174 VSUBS 0.0294f
C5758 VOUT.n1381 VSUBS 0.0689f
C5759 VOUT.n1382 VSUBS 0.03f
C5760 VOUT.n1383 VSUBS 0.0365f
C5761 VOUT.n1384 VSUBS 0.0615f
C5762 VOUT.n1385 VSUBS 0.0195f
C5763 VOUT.n1386 VSUBS 0.00998f
C5764 VOUT.n1387 VSUBS 0.0373f
C5765 VOUT.n1388 VSUBS 0.223f
C5766 VOUT.n1389 VSUBS 0.223f
C5767 VOUT.t304 VSUBS 0.0294f
C5768 VOUT.t310 VSUBS 0.0294f
C5769 VOUT.n1390 VSUBS 0.0689f
C5770 VOUT.n1391 VSUBS 0.03f
C5771 VOUT.n1392 VSUBS 0.0365f
C5772 VOUT.n1393 VSUBS 0.0615f
C5773 VOUT.n1394 VSUBS 0.0195f
C5774 VOUT.n1395 VSUBS 0.00998f
C5775 VOUT.n1396 VSUBS 0.0373f
C5776 VOUT.n1397 VSUBS 0.223f
C5777 VOUT.n1398 VSUBS 0.223f
C5778 VOUT.t232 VSUBS 0.0294f
C5779 VOUT.t152 VSUBS 0.0294f
C5780 VOUT.n1399 VSUBS 0.0689f
C5781 VOUT.n1400 VSUBS 0.03f
C5782 VOUT.n1401 VSUBS 0.0365f
C5783 VOUT.n1402 VSUBS 0.0615f
C5784 VOUT.n1403 VSUBS 0.0195f
C5785 VOUT.n1404 VSUBS 0.00998f
C5786 VOUT.n1405 VSUBS 0.0373f
C5787 VOUT.n1406 VSUBS 0.223f
C5788 VOUT.n1407 VSUBS 0.223f
C5789 VOUT.t194 VSUBS 0.0294f
C5790 VOUT.t295 VSUBS 0.0294f
C5791 VOUT.n1408 VSUBS 0.0689f
C5792 VOUT.n1409 VSUBS 0.03f
C5793 VOUT.n1410 VSUBS 0.0365f
C5794 VOUT.n1411 VSUBS 0.0615f
C5795 VOUT.n1412 VSUBS 0.0195f
C5796 VOUT.n1413 VSUBS 0.00998f
C5797 VOUT.n1414 VSUBS 0.0373f
C5798 VOUT.n1415 VSUBS 0.223f
C5799 VOUT.n1416 VSUBS 0.223f
C5800 VOUT.t277 VSUBS 0.0294f
C5801 VOUT.t186 VSUBS 0.0294f
C5802 VOUT.n1417 VSUBS 0.0689f
C5803 VOUT.n1418 VSUBS 0.03f
C5804 VOUT.n1419 VSUBS 0.0365f
C5805 VOUT.n1420 VSUBS 0.0615f
C5806 VOUT.n1421 VSUBS 0.0195f
C5807 VOUT.n1422 VSUBS 0.00998f
C5808 VOUT.n1423 VSUBS 0.0373f
C5809 VOUT.n1424 VSUBS 0.223f
C5810 VOUT.n1425 VSUBS 0.223f
C5811 VOUT.t172 VSUBS 0.0294f
C5812 VOUT.t328 VSUBS 0.0294f
C5813 VOUT.n1426 VSUBS 0.0689f
C5814 VOUT.n1427 VSUBS 0.03f
C5815 VOUT.n1428 VSUBS 0.0365f
C5816 VOUT.n1429 VSUBS 0.0615f
C5817 VOUT.n1430 VSUBS 0.0195f
C5818 VOUT.n1431 VSUBS 0.00998f
C5819 VOUT.n1432 VSUBS 0.0373f
C5820 VOUT.n1433 VSUBS 0.223f
C5821 VOUT.n1434 VSUBS 0.223f
C5822 VOUT.t233 VSUBS 0.0294f
C5823 VOUT.t299 VSUBS 0.0294f
C5824 VOUT.n1435 VSUBS 0.0689f
C5825 VOUT.n1436 VSUBS 0.03f
C5826 VOUT.n1437 VSUBS 0.0365f
C5827 VOUT.n1438 VSUBS 0.0615f
C5828 VOUT.n1439 VSUBS 0.0195f
C5829 VOUT.n1440 VSUBS 0.00998f
C5830 VOUT.n1441 VSUBS 0.0373f
C5831 VOUT.n1442 VSUBS 0.223f
C5832 VOUT.n1443 VSUBS 0.223f
C5833 VOUT.t305 VSUBS 0.0294f
C5834 VOUT.t154 VSUBS 0.0294f
C5835 VOUT.n1444 VSUBS 0.0689f
C5836 VOUT.n1445 VSUBS 0.03f
C5837 VOUT.n1446 VSUBS 0.0365f
C5838 VOUT.n1447 VSUBS 0.0615f
C5839 VOUT.n1448 VSUBS 0.0195f
C5840 VOUT.n1449 VSUBS 0.00998f
C5841 VOUT.n1450 VSUBS 0.0373f
C5842 VOUT.n1451 VSUBS 0.223f
C5843 VOUT.n1452 VSUBS 0.223f
C5844 VOUT.t167 VSUBS 0.0294f
C5845 VOUT.t250 VSUBS 0.0294f
C5846 VOUT.n1453 VSUBS 0.0689f
C5847 VOUT.n1454 VSUBS 0.03f
C5848 VOUT.n1455 VSUBS 0.0365f
C5849 VOUT.n1456 VSUBS 0.0615f
C5850 VOUT.n1457 VSUBS 0.0195f
C5851 VOUT.n1458 VSUBS 0.00998f
C5852 VOUT.n1459 VSUBS 0.0373f
C5853 VOUT.n1460 VSUBS 0.223f
C5854 VOUT.n1461 VSUBS 0.223f
C5855 VOUT.t279 VSUBS 0.0294f
C5856 VOUT.t177 VSUBS 0.0294f
C5857 VOUT.n1462 VSUBS 0.0689f
C5858 VOUT.n1463 VSUBS 0.03f
C5859 VOUT.n1464 VSUBS 0.0365f
C5860 VOUT.n1465 VSUBS 0.0615f
C5861 VOUT.n1466 VSUBS 0.0195f
C5862 VOUT.n1467 VSUBS 0.00998f
C5863 VOUT.n1468 VSUBS 0.0373f
C5864 VOUT.n1469 VSUBS 0.223f
C5865 VOUT.n1470 VSUBS 0.223f
C5866 VOUT.t146 VSUBS 0.0294f
C5867 VOUT.t228 VSUBS 0.0294f
C5868 VOUT.n1471 VSUBS 0.0689f
C5869 VOUT.n1472 VSUBS 0.03f
C5870 VOUT.n1473 VSUBS 0.0365f
C5871 VOUT.n1474 VSUBS 0.0615f
C5872 VOUT.n1475 VSUBS 0.0195f
C5873 VOUT.n1476 VSUBS 0.00998f
C5874 VOUT.n1477 VSUBS 0.0373f
C5875 VOUT.n1478 VSUBS 0.223f
C5876 VOUT.n1479 VSUBS 0.223f
C5877 VOUT.t307 VSUBS 0.0294f
C5878 VOUT.t296 VSUBS 0.0294f
C5879 VOUT.n1480 VSUBS 0.0689f
C5880 VOUT.n1481 VSUBS 0.03f
C5881 VOUT.n1482 VSUBS 0.0365f
C5882 VOUT.n1483 VSUBS 0.0615f
C5883 VOUT.n1484 VSUBS 0.0195f
C5884 VOUT.n1485 VSUBS 0.00998f
C5885 VOUT.n1486 VSUBS 0.0373f
C5886 VOUT.n1487 VSUBS 0.223f
C5887 VOUT.n1488 VSUBS 0.223f
C5888 VOUT.t297 VSUBS 0.0294f
C5889 VOUT.t208 VSUBS 0.0294f
C5890 VOUT.n1489 VSUBS 0.0689f
C5891 VOUT.n1490 VSUBS 0.03f
C5892 VOUT.n1491 VSUBS 0.0365f
C5893 VOUT.n1492 VSUBS 0.0615f
C5894 VOUT.n1493 VSUBS 0.0195f
C5895 VOUT.n1494 VSUBS 0.00998f
C5896 VOUT.n1495 VSUBS 0.0373f
C5897 VOUT.n1496 VSUBS 0.223f
C5898 VOUT.n1497 VSUBS 0.223f
C5899 VOUT.t199 VSUBS 0.0294f
C5900 VOUT.n1498 VSUBS 0.0982f
C5901 VOUT.n1499 VSUBS 0.03f
C5902 VOUT.n1500 VSUBS 0.0365f
C5903 VOUT.n1501 VSUBS 0.0615f
C5904 VOUT.n1502 VSUBS 0.0195f
C5905 VOUT.n1503 VSUBS 0.00998f
C5906 VOUT.n1504 VSUBS 0.0373f
C5907 VOUT.n1505 VSUBS 0.119f
C5908 VOUT.n1506 VSUBS 0.0358f
C5909 VOUT.n1507 VSUBS 0.041f
C5910 VOUT.n1508 VSUBS 0.0711f
C5911 VOUT.t45 VSUBS 0.0294f
C5912 VOUT.n1509 VSUBS 0.0985f
C5913 VOUT.n1510 VSUBS 0.0181f
C5914 VOUT.n1511 VSUBS 0.00878f
C5915 VOUT.n1512 VSUBS 0.0373f
C5916 VOUT.n1513 VSUBS 0.322f
C5917 VOUT.n1514 VSUBS 0.223f
C5918 VOUT.n1515 VSUBS 0.0358f
C5919 VOUT.n1516 VSUBS 0.0365f
C5920 VOUT.n1517 VSUBS 0.0711f
C5921 VOUT.t369 VSUBS 0.0294f
C5922 VOUT.t357 VSUBS 0.0294f
C5923 VOUT.n1518 VSUBS 0.0691f
C5924 VOUT.n1519 VSUBS 0.0181f
C5925 VOUT.n1520 VSUBS 0.00878f
C5926 VOUT.n1521 VSUBS 0.0373f
C5927 VOUT.n1522 VSUBS 0.223f
C5928 VOUT.n1523 VSUBS 0.223f
C5929 VOUT.n1524 VSUBS 0.0358f
C5930 VOUT.n1525 VSUBS 0.0365f
C5931 VOUT.n1526 VSUBS 0.0711f
C5932 VOUT.t78 VSUBS 0.0294f
C5933 VOUT.t397 VSUBS 0.0294f
C5934 VOUT.n1527 VSUBS 0.0691f
C5935 VOUT.n1528 VSUBS 0.0181f
C5936 VOUT.n1529 VSUBS 0.00878f
C5937 VOUT.n1530 VSUBS 0.0373f
C5938 VOUT.n1531 VSUBS 0.223f
C5939 VOUT.n1532 VSUBS 0.223f
C5940 VOUT.n1533 VSUBS 0.0358f
C5941 VOUT.n1534 VSUBS 0.0365f
C5942 VOUT.n1535 VSUBS 0.0711f
C5943 VOUT.t393 VSUBS 0.0294f
C5944 VOUT.t490 VSUBS 0.0294f
C5945 VOUT.n1536 VSUBS 0.0691f
C5946 VOUT.n1537 VSUBS 0.0181f
C5947 VOUT.n1538 VSUBS 0.00878f
C5948 VOUT.n1539 VSUBS 0.0373f
C5949 VOUT.n1540 VSUBS 0.223f
C5950 VOUT.n1541 VSUBS 0.223f
C5951 VOUT.n1542 VSUBS 0.0358f
C5952 VOUT.n1543 VSUBS 0.0365f
C5953 VOUT.n1544 VSUBS 0.0711f
C5954 VOUT.t52 VSUBS 0.0294f
C5955 VOUT.t355 VSUBS 0.0294f
C5956 VOUT.n1545 VSUBS 0.0691f
C5957 VOUT.n1546 VSUBS 0.0181f
C5958 VOUT.n1547 VSUBS 0.00878f
C5959 VOUT.n1548 VSUBS 0.0373f
C5960 VOUT.n1549 VSUBS 0.223f
C5961 VOUT.n1550 VSUBS 0.223f
C5962 VOUT.n1551 VSUBS 0.0358f
C5963 VOUT.n1552 VSUBS 0.0365f
C5964 VOUT.n1553 VSUBS 0.0711f
C5965 VOUT.t389 VSUBS 0.0294f
C5966 VOUT.t42 VSUBS 0.0294f
C5967 VOUT.n1554 VSUBS 0.0691f
C5968 VOUT.n1555 VSUBS 0.0181f
C5969 VOUT.n1556 VSUBS 0.00878f
C5970 VOUT.n1557 VSUBS 0.0373f
C5971 VOUT.n1558 VSUBS 0.223f
C5972 VOUT.n1559 VSUBS 0.223f
C5973 VOUT.n1560 VSUBS 0.0358f
C5974 VOUT.n1561 VSUBS 0.0365f
C5975 VOUT.n1562 VSUBS 0.0711f
C5976 VOUT.t21 VSUBS 0.0294f
C5977 VOUT.t374 VSUBS 0.0294f
C5978 VOUT.n1563 VSUBS 0.0691f
C5979 VOUT.n1564 VSUBS 0.0181f
C5980 VOUT.n1565 VSUBS 0.00878f
C5981 VOUT.n1566 VSUBS 0.0373f
C5982 VOUT.n1567 VSUBS 0.223f
C5983 VOUT.n1568 VSUBS 0.223f
C5984 VOUT.n1569 VSUBS 0.0358f
C5985 VOUT.n1570 VSUBS 0.0365f
C5986 VOUT.n1571 VSUBS 0.0711f
C5987 VOUT.t430 VSUBS 0.0294f
C5988 VOUT.t512 VSUBS 0.0294f
C5989 VOUT.n1572 VSUBS 0.0691f
C5990 VOUT.n1573 VSUBS 0.0181f
C5991 VOUT.n1574 VSUBS 0.00878f
C5992 VOUT.n1575 VSUBS 0.0373f
C5993 VOUT.n1576 VSUBS 0.223f
C5994 VOUT.n1577 VSUBS 0.223f
C5995 VOUT.n1578 VSUBS 0.0358f
C5996 VOUT.n1579 VSUBS 0.0365f
C5997 VOUT.n1580 VSUBS 0.0711f
C5998 VOUT.t127 VSUBS 0.0294f
C5999 VOUT.t57 VSUBS 0.0294f
C6000 VOUT.n1581 VSUBS 0.0691f
C6001 VOUT.n1582 VSUBS 0.0181f
C6002 VOUT.n1583 VSUBS 0.00878f
C6003 VOUT.n1584 VSUBS 0.0373f
C6004 VOUT.n1585 VSUBS 0.223f
C6005 VOUT.n1586 VSUBS 0.223f
C6006 VOUT.n1587 VSUBS 0.0358f
C6007 VOUT.n1588 VSUBS 0.0365f
C6008 VOUT.n1589 VSUBS 0.0711f
C6009 VOUT.t513 VSUBS 0.0294f
C6010 VOUT.t63 VSUBS 0.0294f
C6011 VOUT.n1590 VSUBS 0.0691f
C6012 VOUT.n1591 VSUBS 0.0181f
C6013 VOUT.n1592 VSUBS 0.00878f
C6014 VOUT.n1593 VSUBS 0.0373f
C6015 VOUT.n1594 VSUBS 0.223f
C6016 VOUT.n1595 VSUBS 0.223f
C6017 VOUT.n1596 VSUBS 0.0358f
C6018 VOUT.n1597 VSUBS 0.0365f
C6019 VOUT.n1598 VSUBS 0.0711f
C6020 VOUT.t134 VSUBS 0.0294f
C6021 VOUT.t17 VSUBS 0.0294f
C6022 VOUT.n1599 VSUBS 0.0691f
C6023 VOUT.n1600 VSUBS 0.0181f
C6024 VOUT.n1601 VSUBS 0.00878f
C6025 VOUT.n1602 VSUBS 0.0373f
C6026 VOUT.n1603 VSUBS 0.223f
C6027 VOUT.n1604 VSUBS 0.223f
C6028 VOUT.n1605 VSUBS 0.0358f
C6029 VOUT.n1606 VSUBS 0.0365f
C6030 VOUT.n1607 VSUBS 0.0711f
C6031 VOUT.t423 VSUBS 0.0294f
C6032 VOUT.t117 VSUBS 0.0294f
C6033 VOUT.n1608 VSUBS 0.0691f
C6034 VOUT.n1609 VSUBS 0.0181f
C6035 VOUT.n1610 VSUBS 0.00878f
C6036 VOUT.n1611 VSUBS 0.0373f
C6037 VOUT.n1612 VSUBS 0.223f
C6038 VOUT.n1613 VSUBS 0.223f
C6039 VOUT.n1614 VSUBS 0.0358f
C6040 VOUT.n1615 VSUBS 0.0365f
C6041 VOUT.n1616 VSUBS 0.0711f
C6042 VOUT.t116 VSUBS 0.0294f
C6043 VOUT.t506 VSUBS 0.0294f
C6044 VOUT.n1617 VSUBS 0.0691f
C6045 VOUT.n1618 VSUBS 0.0181f
C6046 VOUT.n1619 VSUBS 0.00878f
C6047 VOUT.n1620 VSUBS 0.0373f
C6048 VOUT.n1621 VSUBS 0.223f
C6049 VOUT.n1622 VSUBS 0.223f
C6050 VOUT.n1623 VSUBS 0.0358f
C6051 VOUT.n1624 VSUBS 0.0365f
C6052 VOUT.n1625 VSUBS 0.0711f
C6053 VOUT.t104 VSUBS 0.0294f
C6054 VOUT.t418 VSUBS 0.0294f
C6055 VOUT.n1626 VSUBS 0.0691f
C6056 VOUT.n1627 VSUBS 0.0181f
C6057 VOUT.n1628 VSUBS 0.00878f
C6058 VOUT.n1629 VSUBS 0.0373f
C6059 VOUT.n1630 VSUBS 0.223f
C6060 VOUT.n1631 VSUBS 0.223f
C6061 VOUT.n1632 VSUBS 0.0358f
C6062 VOUT.n1633 VSUBS 0.0365f
C6063 VOUT.n1634 VSUBS 0.0711f
C6064 VOUT.t126 VSUBS 0.0294f
C6065 VOUT.t491 VSUBS 0.0294f
C6066 VOUT.n1635 VSUBS 0.0691f
C6067 VOUT.n1636 VSUBS 0.0181f
C6068 VOUT.n1637 VSUBS 0.00878f
C6069 VOUT.n1638 VSUBS 0.0373f
C6070 VOUT.n1639 VSUBS 0.223f
C6071 VOUT.n1640 VSUBS 0.223f
C6072 VOUT.n1641 VSUBS 0.0358f
C6073 VOUT.n1642 VSUBS 0.0365f
C6074 VOUT.n1643 VSUBS 0.0711f
C6075 VOUT.t371 VSUBS 0.0294f
C6076 VOUT.t466 VSUBS 0.0294f
C6077 VOUT.n1644 VSUBS 0.0691f
C6078 VOUT.n1645 VSUBS 0.0181f
C6079 VOUT.n1646 VSUBS 0.00878f
C6080 VOUT.n1647 VSUBS 0.0373f
C6081 VOUT.n1648 VSUBS 0.223f
C6082 VOUT.n1649 VSUBS 0.223f
C6083 VOUT.n1650 VSUBS 0.0358f
C6084 VOUT.n1651 VSUBS 0.0365f
C6085 VOUT.n1652 VSUBS 0.0711f
C6086 VOUT.t377 VSUBS 0.0294f
C6087 VOUT.t64 VSUBS 0.0294f
C6088 VOUT.n1653 VSUBS 0.0691f
C6089 VOUT.n1654 VSUBS 0.0181f
C6090 VOUT.n1655 VSUBS 0.00878f
C6091 VOUT.n1656 VSUBS 0.0373f
C6092 VOUT.n1657 VSUBS 0.223f
C6093 VOUT.n1658 VSUBS 0.223f
C6094 VOUT.n1659 VSUBS 0.0358f
C6095 VOUT.n1660 VSUBS 0.0365f
C6096 VOUT.n1661 VSUBS 0.0711f
C6097 VOUT.t79 VSUBS 0.0294f
C6098 VOUT.t19 VSUBS 0.0294f
C6099 VOUT.n1662 VSUBS 0.0691f
C6100 VOUT.n1663 VSUBS 0.0181f
C6101 VOUT.n1664 VSUBS 0.00878f
C6102 VOUT.n1665 VSUBS 0.0373f
C6103 VOUT.n1666 VSUBS 0.223f
C6104 VOUT.n1667 VSUBS 0.223f
C6105 VOUT.n1668 VSUBS 0.0358f
C6106 VOUT.n1669 VSUBS 0.0365f
C6107 VOUT.n1670 VSUBS 0.0711f
C6108 VOUT.t503 VSUBS 0.0294f
C6109 VOUT.t478 VSUBS 0.0294f
C6110 VOUT.n1671 VSUBS 0.0691f
C6111 VOUT.n1672 VSUBS 0.0181f
C6112 VOUT.n1673 VSUBS 0.00878f
C6113 VOUT.n1674 VSUBS 0.0373f
C6114 VOUT.n1675 VSUBS 0.223f
C6115 VOUT.n1676 VSUBS 0.223f
C6116 VOUT.n1677 VSUBS 0.0358f
C6117 VOUT.n1678 VSUBS 0.0365f
C6118 VOUT.n1679 VSUBS 0.0711f
C6119 VOUT.t406 VSUBS 0.0294f
C6120 VOUT.t132 VSUBS 0.0294f
C6121 VOUT.n1680 VSUBS 0.0691f
C6122 VOUT.n1681 VSUBS 0.0181f
C6123 VOUT.n1682 VSUBS 0.00878f
C6124 VOUT.n1683 VSUBS 0.0373f
C6125 VOUT.n1684 VSUBS 0.223f
C6126 VOUT.n1685 VSUBS 0.223f
C6127 VOUT.n1686 VSUBS 0.0358f
C6128 VOUT.n1687 VSUBS 0.0365f
C6129 VOUT.n1688 VSUBS 0.0711f
C6130 VOUT.t501 VSUBS 0.0294f
C6131 VOUT.n1689 VSUBS 0.0985f
C6132 VOUT.n1690 VSUBS 0.0181f
C6133 VOUT.n1691 VSUBS 0.00878f
C6134 VOUT.n1692 VSUBS 0.0373f
C6135 VOUT.n1693 VSUBS 0.119f
C6136 VOUT.t22 VSUBS 0.0294f
C6137 VOUT.n1694 VSUBS 0.0984f
C6138 VOUT.n1695 VSUBS 0.0316f
C6139 VOUT.n1696 VSUBS 0.041f
C6140 VOUT.n1697 VSUBS 0.0655f
C6141 VOUT.n1698 VSUBS 0.019f
C6142 VOUT.n1699 VSUBS 0.0094f
C6143 VOUT.n1700 VSUBS 0.0373f
C6144 VOUT.n1701 VSUBS 0.322f
C6145 VOUT.n1702 VSUBS 0.223f
C6146 VOUT.t422 VSUBS 0.0294f
C6147 VOUT.t105 VSUBS 0.0294f
C6148 VOUT.n1703 VSUBS 0.069f
C6149 VOUT.n1704 VSUBS 0.0316f
C6150 VOUT.n1705 VSUBS 0.0365f
C6151 VOUT.n1706 VSUBS 0.0655f
C6152 VOUT.n1707 VSUBS 0.019f
C6153 VOUT.n1708 VSUBS 0.0094f
C6154 VOUT.n1709 VSUBS 0.0373f
C6155 VOUT.n1710 VSUBS 0.223f
C6156 VOUT.n1711 VSUBS 0.223f
C6157 VOUT.t130 VSUBS 0.0294f
C6158 VOUT.t62 VSUBS 0.0294f
C6159 VOUT.n1712 VSUBS 0.069f
C6160 VOUT.n1713 VSUBS 0.0316f
C6161 VOUT.n1714 VSUBS 0.0365f
C6162 VOUT.n1715 VSUBS 0.0655f
C6163 VOUT.n1716 VSUBS 0.019f
C6164 VOUT.n1717 VSUBS 0.0094f
C6165 VOUT.n1718 VSUBS 0.0373f
C6166 VOUT.n1719 VSUBS 0.223f
C6167 VOUT.n1720 VSUBS 0.223f
C6168 VOUT.t404 VSUBS 0.0294f
C6169 VOUT.t66 VSUBS 0.0294f
C6170 VOUT.n1721 VSUBS 0.069f
C6171 VOUT.n1722 VSUBS 0.0316f
C6172 VOUT.n1723 VSUBS 0.0365f
C6173 VOUT.n1724 VSUBS 0.0655f
C6174 VOUT.n1725 VSUBS 0.019f
C6175 VOUT.n1726 VSUBS 0.0094f
C6176 VOUT.n1727 VSUBS 0.0373f
C6177 VOUT.n1728 VSUBS 0.223f
C6178 VOUT.n1729 VSUBS 0.223f
C6179 VOUT.t412 VSUBS 0.0294f
C6180 VOUT.t59 VSUBS 0.0294f
C6181 VOUT.n1730 VSUBS 0.069f
C6182 VOUT.n1731 VSUBS 0.0316f
C6183 VOUT.n1732 VSUBS 0.0365f
C6184 VOUT.n1733 VSUBS 0.0655f
C6185 VOUT.n1734 VSUBS 0.019f
C6186 VOUT.n1735 VSUBS 0.0094f
C6187 VOUT.n1736 VSUBS 0.0373f
C6188 VOUT.n1737 VSUBS 0.223f
C6189 VOUT.n1738 VSUBS 0.223f
C6190 VOUT.t76 VSUBS 0.0294f
C6191 VOUT.t88 VSUBS 0.0294f
C6192 VOUT.n1739 VSUBS 0.069f
C6193 VOUT.n1740 VSUBS 0.0316f
C6194 VOUT.n1741 VSUBS 0.0365f
C6195 VOUT.n1742 VSUBS 0.0655f
C6196 VOUT.n1743 VSUBS 0.019f
C6197 VOUT.n1744 VSUBS 0.0094f
C6198 VOUT.n1745 VSUBS 0.0373f
C6199 VOUT.n1746 VSUBS 0.223f
C6200 VOUT.n1747 VSUBS 0.223f
C6201 VOUT.t75 VSUBS 0.0294f
C6202 VOUT.t379 VSUBS 0.0294f
C6203 VOUT.n1748 VSUBS 0.069f
C6204 VOUT.n1749 VSUBS 0.0316f
C6205 VOUT.n1750 VSUBS 0.0365f
C6206 VOUT.n1751 VSUBS 0.0655f
C6207 VOUT.n1752 VSUBS 0.019f
C6208 VOUT.n1753 VSUBS 0.0094f
C6209 VOUT.n1754 VSUBS 0.0373f
C6210 VOUT.n1755 VSUBS 0.223f
C6211 VOUT.n1756 VSUBS 0.223f
C6212 VOUT.t441 VSUBS 0.0294f
C6213 VOUT.t375 VSUBS 0.0294f
C6214 VOUT.n1757 VSUBS 0.069f
C6215 VOUT.n1758 VSUBS 0.0316f
C6216 VOUT.n1759 VSUBS 0.0365f
C6217 VOUT.n1760 VSUBS 0.0655f
C6218 VOUT.n1761 VSUBS 0.019f
C6219 VOUT.n1762 VSUBS 0.0094f
C6220 VOUT.n1763 VSUBS 0.0373f
C6221 VOUT.n1764 VSUBS 0.223f
C6222 VOUT.n1765 VSUBS 0.223f
C6223 VOUT.t24 VSUBS 0.0294f
C6224 VOUT.t61 VSUBS 0.0294f
C6225 VOUT.n1766 VSUBS 0.069f
C6226 VOUT.n1767 VSUBS 0.0316f
C6227 VOUT.n1768 VSUBS 0.0365f
C6228 VOUT.n1769 VSUBS 0.0655f
C6229 VOUT.n1770 VSUBS 0.019f
C6230 VOUT.n1771 VSUBS 0.0094f
C6231 VOUT.n1772 VSUBS 0.0373f
C6232 VOUT.n1773 VSUBS 0.223f
C6233 VOUT.n1774 VSUBS 0.223f
C6234 VOUT.t414 VSUBS 0.0294f
C6235 VOUT.t500 VSUBS 0.0294f
C6236 VOUT.n1775 VSUBS 0.069f
C6237 VOUT.n1776 VSUBS 0.0316f
C6238 VOUT.n1777 VSUBS 0.0365f
C6239 VOUT.n1778 VSUBS 0.0655f
C6240 VOUT.n1779 VSUBS 0.019f
C6241 VOUT.n1780 VSUBS 0.0094f
C6242 VOUT.n1781 VSUBS 0.0373f
C6243 VOUT.n1782 VSUBS 0.223f
C6244 VOUT.n1783 VSUBS 0.223f
C6245 VOUT.t351 VSUBS 0.0294f
C6246 VOUT.t23 VSUBS 0.0294f
C6247 VOUT.n1784 VSUBS 0.069f
C6248 VOUT.n1785 VSUBS 0.0316f
C6249 VOUT.n1786 VSUBS 0.0365f
C6250 VOUT.n1787 VSUBS 0.0655f
C6251 VOUT.n1788 VSUBS 0.019f
C6252 VOUT.n1789 VSUBS 0.0094f
C6253 VOUT.n1790 VSUBS 0.0373f
C6254 VOUT.n1791 VSUBS 0.223f
C6255 VOUT.n1792 VSUBS 0.223f
C6256 VOUT.t342 VSUBS 0.0294f
C6257 VOUT.t27 VSUBS 0.0294f
C6258 VOUT.n1793 VSUBS 0.069f
C6259 VOUT.n1794 VSUBS 0.0316f
C6260 VOUT.n1795 VSUBS 0.0365f
C6261 VOUT.n1796 VSUBS 0.0655f
C6262 VOUT.n1797 VSUBS 0.019f
C6263 VOUT.n1798 VSUBS 0.0094f
C6264 VOUT.n1799 VSUBS 0.0373f
C6265 VOUT.n1800 VSUBS 0.223f
C6266 VOUT.n1801 VSUBS 0.223f
C6267 VOUT.t40 VSUBS 0.0294f
C6268 VOUT.t497 VSUBS 0.0294f
C6269 VOUT.n1802 VSUBS 0.069f
C6270 VOUT.n1803 VSUBS 0.0316f
C6271 VOUT.n1804 VSUBS 0.0365f
C6272 VOUT.n1805 VSUBS 0.0655f
C6273 VOUT.n1806 VSUBS 0.019f
C6274 VOUT.n1807 VSUBS 0.0094f
C6275 VOUT.n1808 VSUBS 0.0373f
C6276 VOUT.n1809 VSUBS 0.223f
C6277 VOUT.n1810 VSUBS 0.223f
C6278 VOUT.t13 VSUBS 0.0294f
C6279 VOUT.t388 VSUBS 0.0294f
C6280 VOUT.n1811 VSUBS 0.069f
C6281 VOUT.n1812 VSUBS 0.0316f
C6282 VOUT.n1813 VSUBS 0.0365f
C6283 VOUT.n1814 VSUBS 0.0655f
C6284 VOUT.n1815 VSUBS 0.019f
C6285 VOUT.n1816 VSUBS 0.0094f
C6286 VOUT.n1817 VSUBS 0.0373f
C6287 VOUT.n1818 VSUBS 0.223f
C6288 VOUT.n1819 VSUBS 0.223f
C6289 VOUT.t114 VSUBS 0.0294f
C6290 VOUT.t73 VSUBS 0.0294f
C6291 VOUT.n1820 VSUBS 0.069f
C6292 VOUT.n1821 VSUBS 0.0316f
C6293 VOUT.n1822 VSUBS 0.0365f
C6294 VOUT.n1823 VSUBS 0.0655f
C6295 VOUT.n1824 VSUBS 0.019f
C6296 VOUT.n1825 VSUBS 0.0094f
C6297 VOUT.n1826 VSUBS 0.0373f
C6298 VOUT.n1827 VSUBS 0.223f
C6299 VOUT.n1828 VSUBS 0.223f
C6300 VOUT.t5 VSUBS 0.0294f
C6301 VOUT.t29 VSUBS 0.0294f
C6302 VOUT.n1829 VSUBS 0.069f
C6303 VOUT.n1830 VSUBS 0.0316f
C6304 VOUT.n1831 VSUBS 0.0365f
C6305 VOUT.n1832 VSUBS 0.0655f
C6306 VOUT.n1833 VSUBS 0.019f
C6307 VOUT.n1834 VSUBS 0.0094f
C6308 VOUT.n1835 VSUBS 0.0373f
C6309 VOUT.n1836 VSUBS 0.223f
C6310 VOUT.n1837 VSUBS 0.223f
C6311 VOUT.t118 VSUBS 0.0294f
C6312 VOUT.t68 VSUBS 0.0294f
C6313 VOUT.n1838 VSUBS 0.069f
C6314 VOUT.n1839 VSUBS 0.0316f
C6315 VOUT.n1840 VSUBS 0.0365f
C6316 VOUT.n1841 VSUBS 0.0655f
C6317 VOUT.n1842 VSUBS 0.019f
C6318 VOUT.n1843 VSUBS 0.0094f
C6319 VOUT.n1844 VSUBS 0.0373f
C6320 VOUT.n1845 VSUBS 0.223f
C6321 VOUT.n1846 VSUBS 0.223f
C6322 VOUT.t489 VSUBS 0.0294f
C6323 VOUT.t427 VSUBS 0.0294f
C6324 VOUT.n1847 VSUBS 0.069f
C6325 VOUT.n1848 VSUBS 0.0316f
C6326 VOUT.n1849 VSUBS 0.0365f
C6327 VOUT.n1850 VSUBS 0.0655f
C6328 VOUT.n1851 VSUBS 0.019f
C6329 VOUT.n1852 VSUBS 0.0094f
C6330 VOUT.n1853 VSUBS 0.0373f
C6331 VOUT.n1854 VSUBS 0.223f
C6332 VOUT.n1855 VSUBS 0.223f
C6333 VOUT.t120 VSUBS 0.0294f
C6334 VOUT.t366 VSUBS 0.0294f
C6335 VOUT.n1856 VSUBS 0.069f
C6336 VOUT.n1857 VSUBS 0.0316f
C6337 VOUT.n1858 VSUBS 0.0365f
C6338 VOUT.n1859 VSUBS 0.0655f
C6339 VOUT.n1860 VSUBS 0.019f
C6340 VOUT.n1861 VSUBS 0.0094f
C6341 VOUT.n1862 VSUBS 0.0373f
C6342 VOUT.n1863 VSUBS 0.223f
C6343 VOUT.n1864 VSUBS 0.223f
C6344 VOUT.t487 VSUBS 0.0294f
C6345 VOUT.t34 VSUBS 0.0294f
C6346 VOUT.n1865 VSUBS 0.069f
C6347 VOUT.n1866 VSUBS 0.0316f
C6348 VOUT.n1867 VSUBS 0.0365f
C6349 VOUT.n1868 VSUBS 0.0655f
C6350 VOUT.n1869 VSUBS 0.019f
C6351 VOUT.n1870 VSUBS 0.0094f
C6352 VOUT.n1871 VSUBS 0.0373f
C6353 VOUT.n1872 VSUBS 0.223f
C6354 VOUT.n1873 VSUBS 0.223f
C6355 VOUT.t440 VSUBS 0.0294f
C6356 VOUT.n1874 VSUBS 0.0984f
C6357 VOUT.n1875 VSUBS 0.0316f
C6358 VOUT.n1876 VSUBS 0.0365f
C6359 VOUT.n1877 VSUBS 0.0655f
C6360 VOUT.n1878 VSUBS 0.019f
C6361 VOUT.n1879 VSUBS 0.0094f
C6362 VOUT.n1880 VSUBS 0.0373f
C6363 VOUT.n1881 VSUBS 0.119f
C6364 VOUT.t87 VSUBS 0.0294f
C6365 VOUT.n1882 VSUBS 0.0983f
C6366 VOUT.n1883 VSUBS 0.0312f
C6367 VOUT.n1884 VSUBS 0.041f
C6368 VOUT.n1885 VSUBS 0.0646f
C6369 VOUT.n1886 VSUBS 0.0191f
C6370 VOUT.n1887 VSUBS 0.00957f
C6371 VOUT.n1888 VSUBS 0.0373f
C6372 VOUT.n1889 VSUBS 0.322f
C6373 VOUT.n1890 VSUBS 0.223f
C6374 VOUT.t95 VSUBS 0.0294f
C6375 VOUT.t488 VSUBS 0.0294f
C6376 VOUT.n1891 VSUBS 0.069f
C6377 VOUT.n1892 VSUBS 0.0312f
C6378 VOUT.n1893 VSUBS 0.0365f
C6379 VOUT.n1894 VSUBS 0.0646f
C6380 VOUT.n1895 VSUBS 0.0191f
C6381 VOUT.n1896 VSUBS 0.00957f
C6382 VOUT.n1897 VSUBS 0.0373f
C6383 VOUT.n1898 VSUBS 0.223f
C6384 VOUT.n1899 VSUBS 0.223f
C6385 VOUT.t361 VSUBS 0.0294f
C6386 VOUT.t415 VSUBS 0.0294f
C6387 VOUT.n1900 VSUBS 0.069f
C6388 VOUT.n1901 VSUBS 0.0312f
C6389 VOUT.n1902 VSUBS 0.0365f
C6390 VOUT.n1903 VSUBS 0.0646f
C6391 VOUT.n1904 VSUBS 0.0191f
C6392 VOUT.n1905 VSUBS 0.00957f
C6393 VOUT.n1906 VSUBS 0.0373f
C6394 VOUT.n1907 VSUBS 0.223f
C6395 VOUT.n1908 VSUBS 0.223f
C6396 VOUT.t368 VSUBS 0.0294f
C6397 VOUT.t131 VSUBS 0.0294f
C6398 VOUT.n1909 VSUBS 0.069f
C6399 VOUT.n1910 VSUBS 0.0312f
C6400 VOUT.n1911 VSUBS 0.0365f
C6401 VOUT.n1912 VSUBS 0.0646f
C6402 VOUT.n1913 VSUBS 0.0191f
C6403 VOUT.n1914 VSUBS 0.00957f
C6404 VOUT.n1915 VSUBS 0.0373f
C6405 VOUT.n1916 VSUBS 0.223f
C6406 VOUT.n1917 VSUBS 0.223f
C6407 VOUT.t91 VSUBS 0.0294f
C6408 VOUT.t390 VSUBS 0.0294f
C6409 VOUT.n1918 VSUBS 0.069f
C6410 VOUT.n1919 VSUBS 0.0312f
C6411 VOUT.n1920 VSUBS 0.0365f
C6412 VOUT.n1921 VSUBS 0.0646f
C6413 VOUT.n1922 VSUBS 0.0191f
C6414 VOUT.n1923 VSUBS 0.00957f
C6415 VOUT.n1924 VSUBS 0.0373f
C6416 VOUT.n1925 VSUBS 0.223f
C6417 VOUT.n1926 VSUBS 0.223f
C6418 VOUT.t93 VSUBS 0.0294f
C6419 VOUT.t483 VSUBS 0.0294f
C6420 VOUT.n1927 VSUBS 0.069f
C6421 VOUT.n1928 VSUBS 0.0312f
C6422 VOUT.n1929 VSUBS 0.0365f
C6423 VOUT.n1930 VSUBS 0.0646f
C6424 VOUT.n1931 VSUBS 0.0191f
C6425 VOUT.n1932 VSUBS 0.00957f
C6426 VOUT.n1933 VSUBS 0.0373f
C6427 VOUT.n1934 VSUBS 0.223f
C6428 VOUT.n1935 VSUBS 0.223f
C6429 VOUT.t122 VSUBS 0.0294f
C6430 VOUT.t94 VSUBS 0.0294f
C6431 VOUT.n1936 VSUBS 0.069f
C6432 VOUT.n1937 VSUBS 0.0312f
C6433 VOUT.n1938 VSUBS 0.0365f
C6434 VOUT.n1939 VSUBS 0.0646f
C6435 VOUT.n1940 VSUBS 0.0191f
C6436 VOUT.n1941 VSUBS 0.00957f
C6437 VOUT.n1942 VSUBS 0.0373f
C6438 VOUT.n1943 VSUBS 0.223f
C6439 VOUT.n1944 VSUBS 0.223f
C6440 VOUT.t100 VSUBS 0.0294f
C6441 VOUT.t48 VSUBS 0.0294f
C6442 VOUT.n1945 VSUBS 0.069f
C6443 VOUT.n1946 VSUBS 0.0312f
C6444 VOUT.n1947 VSUBS 0.0365f
C6445 VOUT.n1948 VSUBS 0.0646f
C6446 VOUT.n1949 VSUBS 0.0191f
C6447 VOUT.n1950 VSUBS 0.00957f
C6448 VOUT.n1951 VSUBS 0.0373f
C6449 VOUT.n1952 VSUBS 0.223f
C6450 VOUT.n1953 VSUBS 0.223f
C6451 VOUT.t394 VSUBS 0.0294f
C6452 VOUT.t464 VSUBS 0.0294f
C6453 VOUT.n1954 VSUBS 0.069f
C6454 VOUT.n1955 VSUBS 0.0312f
C6455 VOUT.n1956 VSUBS 0.0365f
C6456 VOUT.n1957 VSUBS 0.0646f
C6457 VOUT.n1958 VSUBS 0.0191f
C6458 VOUT.n1959 VSUBS 0.00957f
C6459 VOUT.n1960 VSUBS 0.0373f
C6460 VOUT.n1961 VSUBS 0.223f
C6461 VOUT.n1962 VSUBS 0.223f
C6462 VOUT.t106 VSUBS 0.0294f
C6463 VOUT.t81 VSUBS 0.0294f
C6464 VOUT.n1963 VSUBS 0.069f
C6465 VOUT.n1964 VSUBS 0.0312f
C6466 VOUT.n1965 VSUBS 0.0365f
C6467 VOUT.n1966 VSUBS 0.0646f
C6468 VOUT.n1967 VSUBS 0.0191f
C6469 VOUT.n1968 VSUBS 0.00957f
C6470 VOUT.n1969 VSUBS 0.0373f
C6471 VOUT.n1970 VSUBS 0.223f
C6472 VOUT.n1971 VSUBS 0.223f
C6473 VOUT.t121 VSUBS 0.0294f
C6474 VOUT.t413 VSUBS 0.0294f
C6475 VOUT.n1972 VSUBS 0.069f
C6476 VOUT.n1973 VSUBS 0.0312f
C6477 VOUT.n1974 VSUBS 0.0365f
C6478 VOUT.n1975 VSUBS 0.0646f
C6479 VOUT.n1976 VSUBS 0.0191f
C6480 VOUT.n1977 VSUBS 0.00957f
C6481 VOUT.n1978 VSUBS 0.0373f
C6482 VOUT.n1979 VSUBS 0.223f
C6483 VOUT.n1980 VSUBS 0.223f
C6484 VOUT.t421 VSUBS 0.0294f
C6485 VOUT.t96 VSUBS 0.0294f
C6486 VOUT.n1981 VSUBS 0.069f
C6487 VOUT.n1982 VSUBS 0.0312f
C6488 VOUT.n1983 VSUBS 0.0365f
C6489 VOUT.n1984 VSUBS 0.0646f
C6490 VOUT.n1985 VSUBS 0.0191f
C6491 VOUT.n1986 VSUBS 0.00957f
C6492 VOUT.n1987 VSUBS 0.0373f
C6493 VOUT.n1988 VSUBS 0.223f
C6494 VOUT.n1989 VSUBS 0.223f
C6495 VOUT.t47 VSUBS 0.0294f
C6496 VOUT.t492 VSUBS 0.0294f
C6497 VOUT.n1990 VSUBS 0.069f
C6498 VOUT.n1991 VSUBS 0.0312f
C6499 VOUT.n1992 VSUBS 0.0365f
C6500 VOUT.n1993 VSUBS 0.0646f
C6501 VOUT.n1994 VSUBS 0.0191f
C6502 VOUT.n1995 VSUBS 0.00957f
C6503 VOUT.n1996 VSUBS 0.0373f
C6504 VOUT.n1997 VSUBS 0.223f
C6505 VOUT.n1998 VSUBS 0.223f
C6506 VOUT.t103 VSUBS 0.0294f
C6507 VOUT.t350 VSUBS 0.0294f
C6508 VOUT.n1999 VSUBS 0.069f
C6509 VOUT.n2000 VSUBS 0.0312f
C6510 VOUT.n2001 VSUBS 0.0365f
C6511 VOUT.n2002 VSUBS 0.0646f
C6512 VOUT.n2003 VSUBS 0.0191f
C6513 VOUT.n2004 VSUBS 0.00957f
C6514 VOUT.n2005 VSUBS 0.0373f
C6515 VOUT.n2006 VSUBS 0.223f
C6516 VOUT.n2007 VSUBS 0.223f
C6517 VOUT.t438 VSUBS 0.0294f
C6518 VOUT.t92 VSUBS 0.0294f
C6519 VOUT.n2008 VSUBS 0.069f
C6520 VOUT.n2009 VSUBS 0.0312f
C6521 VOUT.n2010 VSUBS 0.0365f
C6522 VOUT.n2011 VSUBS 0.0646f
C6523 VOUT.n2012 VSUBS 0.0191f
C6524 VOUT.n2013 VSUBS 0.00957f
C6525 VOUT.n2014 VSUBS 0.0373f
C6526 VOUT.n2015 VSUBS 0.223f
C6527 VOUT.n2016 VSUBS 0.223f
C6528 VOUT.t46 VSUBS 0.0294f
C6529 VOUT.t51 VSUBS 0.0294f
C6530 VOUT.n2017 VSUBS 0.069f
C6531 VOUT.n2018 VSUBS 0.0312f
C6532 VOUT.n2019 VSUBS 0.0365f
C6533 VOUT.n2020 VSUBS 0.0646f
C6534 VOUT.n2021 VSUBS 0.0191f
C6535 VOUT.n2022 VSUBS 0.00957f
C6536 VOUT.n2023 VSUBS 0.0373f
C6537 VOUT.n2024 VSUBS 0.223f
C6538 VOUT.n2025 VSUBS 0.223f
C6539 VOUT.t391 VSUBS 0.0294f
C6540 VOUT.t384 VSUBS 0.0294f
C6541 VOUT.n2026 VSUBS 0.069f
C6542 VOUT.n2027 VSUBS 0.0312f
C6543 VOUT.n2028 VSUBS 0.0365f
C6544 VOUT.n2029 VSUBS 0.0646f
C6545 VOUT.n2030 VSUBS 0.0191f
C6546 VOUT.n2031 VSUBS 0.00957f
C6547 VOUT.n2032 VSUBS 0.0373f
C6548 VOUT.n2033 VSUBS 0.223f
C6549 VOUT.n2034 VSUBS 0.223f
C6550 VOUT.t25 VSUBS 0.0294f
C6551 VOUT.t349 VSUBS 0.0294f
C6552 VOUT.n2035 VSUBS 0.069f
C6553 VOUT.n2036 VSUBS 0.0312f
C6554 VOUT.n2037 VSUBS 0.0365f
C6555 VOUT.n2038 VSUBS 0.0646f
C6556 VOUT.n2039 VSUBS 0.0191f
C6557 VOUT.n2040 VSUBS 0.00957f
C6558 VOUT.n2041 VSUBS 0.0373f
C6559 VOUT.n2042 VSUBS 0.223f
C6560 VOUT.n2043 VSUBS 0.223f
C6561 VOUT.t37 VSUBS 0.0294f
C6562 VOUT.t109 VSUBS 0.0294f
C6563 VOUT.n2044 VSUBS 0.069f
C6564 VOUT.n2045 VSUBS 0.0312f
C6565 VOUT.n2046 VSUBS 0.0365f
C6566 VOUT.n2047 VSUBS 0.0646f
C6567 VOUT.n2048 VSUBS 0.0191f
C6568 VOUT.n2049 VSUBS 0.00957f
C6569 VOUT.n2050 VSUBS 0.0373f
C6570 VOUT.n2051 VSUBS 0.223f
C6571 VOUT.n2052 VSUBS 0.223f
C6572 VOUT.t494 VSUBS 0.0294f
C6573 VOUT.t386 VSUBS 0.0294f
C6574 VOUT.n2053 VSUBS 0.069f
C6575 VOUT.n2054 VSUBS 0.0312f
C6576 VOUT.n2055 VSUBS 0.0365f
C6577 VOUT.n2056 VSUBS 0.0646f
C6578 VOUT.n2057 VSUBS 0.0191f
C6579 VOUT.n2058 VSUBS 0.00957f
C6580 VOUT.n2059 VSUBS 0.0373f
C6581 VOUT.n2060 VSUBS 0.223f
C6582 VOUT.n2061 VSUBS 0.223f
C6583 VOUT.t385 VSUBS 0.0294f
C6584 VOUT.n2062 VSUBS 0.0983f
C6585 VOUT.n2063 VSUBS 0.0312f
C6586 VOUT.n2064 VSUBS 0.0365f
C6587 VOUT.n2065 VSUBS 0.0646f
C6588 VOUT.n2066 VSUBS 0.0191f
C6589 VOUT.n2067 VSUBS 0.00957f
C6590 VOUT.n2068 VSUBS 0.0373f
C6591 VOUT.n2069 VSUBS 0.119f
C6592 VOUT.t26 VSUBS 0.0294f
C6593 VOUT.n2070 VSUBS 0.0984f
C6594 VOUT.n2071 VSUBS 0.0324f
C6595 VOUT.n2072 VSUBS 0.041f
C6596 VOUT.n2073 VSUBS 0.0678f
C6597 VOUT.n2074 VSUBS 0.0188f
C6598 VOUT.n2075 VSUBS 0.00925f
C6599 VOUT.n2076 VSUBS 0.0373f
C6600 VOUT.n2077 VSUBS 0.322f
C6601 VOUT.n2078 VSUBS 0.223f
C6602 VOUT.t102 VSUBS 0.0294f
C6603 VOUT.t493 VSUBS 0.0294f
C6604 VOUT.n2079 VSUBS 0.069f
C6605 VOUT.n2080 VSUBS 0.0324f
C6606 VOUT.n2081 VSUBS 0.0365f
C6607 VOUT.n2082 VSUBS 0.0678f
C6608 VOUT.n2083 VSUBS 0.0188f
C6609 VOUT.n2084 VSUBS 0.00925f
C6610 VOUT.n2085 VSUBS 0.0373f
C6611 VOUT.n2086 VSUBS 0.223f
C6612 VOUT.n2087 VSUBS 0.223f
C6613 VOUT.t502 VSUBS 0.0294f
C6614 VOUT.t372 VSUBS 0.0294f
C6615 VOUT.n2088 VSUBS 0.069f
C6616 VOUT.n2089 VSUBS 0.0324f
C6617 VOUT.n2090 VSUBS 0.0365f
C6618 VOUT.n2091 VSUBS 0.0678f
C6619 VOUT.n2092 VSUBS 0.0188f
C6620 VOUT.n2093 VSUBS 0.00925f
C6621 VOUT.n2094 VSUBS 0.0373f
C6622 VOUT.n2095 VSUBS 0.223f
C6623 VOUT.n2096 VSUBS 0.223f
C6624 VOUT.t419 VSUBS 0.0294f
C6625 VOUT.t485 VSUBS 0.0294f
C6626 VOUT.n2097 VSUBS 0.069f
C6627 VOUT.n2098 VSUBS 0.0324f
C6628 VOUT.n2099 VSUBS 0.0365f
C6629 VOUT.n2100 VSUBS 0.0678f
C6630 VOUT.n2101 VSUBS 0.0188f
C6631 VOUT.n2102 VSUBS 0.00925f
C6632 VOUT.n2103 VSUBS 0.0373f
C6633 VOUT.n2104 VSUBS 0.223f
C6634 VOUT.n2105 VSUBS 0.223f
C6635 VOUT.t428 VSUBS 0.0294f
C6636 VOUT.t499 VSUBS 0.0294f
C6637 VOUT.n2106 VSUBS 0.069f
C6638 VOUT.n2107 VSUBS 0.0324f
C6639 VOUT.n2108 VSUBS 0.0365f
C6640 VOUT.n2109 VSUBS 0.0678f
C6641 VOUT.n2110 VSUBS 0.0188f
C6642 VOUT.n2111 VSUBS 0.00925f
C6643 VOUT.n2112 VSUBS 0.0373f
C6644 VOUT.n2113 VSUBS 0.223f
C6645 VOUT.n2114 VSUBS 0.223f
C6646 VOUT.t74 VSUBS 0.0294f
C6647 VOUT.t356 VSUBS 0.0294f
C6648 VOUT.n2115 VSUBS 0.069f
C6649 VOUT.n2116 VSUBS 0.0324f
C6650 VOUT.n2117 VSUBS 0.0365f
C6651 VOUT.n2118 VSUBS 0.0678f
C6652 VOUT.n2119 VSUBS 0.0188f
C6653 VOUT.n2120 VSUBS 0.00925f
C6654 VOUT.n2121 VSUBS 0.0373f
C6655 VOUT.n2122 VSUBS 0.223f
C6656 VOUT.n2123 VSUBS 0.223f
C6657 VOUT.t429 VSUBS 0.0294f
C6658 VOUT.t353 VSUBS 0.0294f
C6659 VOUT.n2124 VSUBS 0.069f
C6660 VOUT.n2125 VSUBS 0.0324f
C6661 VOUT.n2126 VSUBS 0.0365f
C6662 VOUT.n2127 VSUBS 0.0678f
C6663 VOUT.n2128 VSUBS 0.0188f
C6664 VOUT.n2129 VSUBS 0.00925f
C6665 VOUT.n2130 VSUBS 0.0373f
C6666 VOUT.n2131 VSUBS 0.223f
C6667 VOUT.n2132 VSUBS 0.223f
C6668 VOUT.t90 VSUBS 0.0294f
C6669 VOUT.t41 VSUBS 0.0294f
C6670 VOUT.n2133 VSUBS 0.069f
C6671 VOUT.n2134 VSUBS 0.0324f
C6672 VOUT.n2135 VSUBS 0.0365f
C6673 VOUT.n2136 VSUBS 0.0678f
C6674 VOUT.n2137 VSUBS 0.0188f
C6675 VOUT.n2138 VSUBS 0.00925f
C6676 VOUT.n2139 VSUBS 0.0373f
C6677 VOUT.n2140 VSUBS 0.223f
C6678 VOUT.n2141 VSUBS 0.223f
C6679 VOUT.t72 VSUBS 0.0294f
C6680 VOUT.t370 VSUBS 0.0294f
C6681 VOUT.n2142 VSUBS 0.069f
C6682 VOUT.n2143 VSUBS 0.0324f
C6683 VOUT.n2144 VSUBS 0.0365f
C6684 VOUT.n2145 VSUBS 0.0678f
C6685 VOUT.n2146 VSUBS 0.0188f
C6686 VOUT.n2147 VSUBS 0.00925f
C6687 VOUT.n2148 VSUBS 0.0373f
C6688 VOUT.n2149 VSUBS 0.223f
C6689 VOUT.n2150 VSUBS 0.223f
C6690 VOUT.t129 VSUBS 0.0294f
C6691 VOUT.t67 VSUBS 0.0294f
C6692 VOUT.n2151 VSUBS 0.069f
C6693 VOUT.n2152 VSUBS 0.0324f
C6694 VOUT.n2153 VSUBS 0.0365f
C6695 VOUT.n2154 VSUBS 0.0678f
C6696 VOUT.n2155 VSUBS 0.0188f
C6697 VOUT.n2156 VSUBS 0.00925f
C6698 VOUT.n2157 VSUBS 0.0373f
C6699 VOUT.n2158 VSUBS 0.223f
C6700 VOUT.n2159 VSUBS 0.223f
C6701 VOUT.t85 VSUBS 0.0294f
C6702 VOUT.t119 VSUBS 0.0294f
C6703 VOUT.n2160 VSUBS 0.069f
C6704 VOUT.n2161 VSUBS 0.0324f
C6705 VOUT.n2162 VSUBS 0.0365f
C6706 VOUT.n2163 VSUBS 0.0678f
C6707 VOUT.n2164 VSUBS 0.0188f
C6708 VOUT.n2165 VSUBS 0.00925f
C6709 VOUT.n2166 VSUBS 0.0373f
C6710 VOUT.n2167 VSUBS 0.223f
C6711 VOUT.n2168 VSUBS 0.223f
C6712 VOUT.t110 VSUBS 0.0294f
C6713 VOUT.t56 VSUBS 0.0294f
C6714 VOUT.n2169 VSUBS 0.069f
C6715 VOUT.n2170 VSUBS 0.0324f
C6716 VOUT.n2171 VSUBS 0.0365f
C6717 VOUT.n2172 VSUBS 0.0678f
C6718 VOUT.n2173 VSUBS 0.0188f
C6719 VOUT.n2174 VSUBS 0.00925f
C6720 VOUT.n2175 VSUBS 0.0373f
C6721 VOUT.n2176 VSUBS 0.223f
C6722 VOUT.n2177 VSUBS 0.223f
C6723 VOUT.t463 VSUBS 0.0294f
C6724 VOUT.t124 VSUBS 0.0294f
C6725 VOUT.n2178 VSUBS 0.069f
C6726 VOUT.n2179 VSUBS 0.0324f
C6727 VOUT.n2180 VSUBS 0.0365f
C6728 VOUT.n2181 VSUBS 0.0678f
C6729 VOUT.n2182 VSUBS 0.0188f
C6730 VOUT.n2183 VSUBS 0.00925f
C6731 VOUT.n2184 VSUBS 0.0373f
C6732 VOUT.n2185 VSUBS 0.223f
C6733 VOUT.n2186 VSUBS 0.223f
C6734 VOUT.t395 VSUBS 0.0294f
C6735 VOUT.t486 VSUBS 0.0294f
C6736 VOUT.n2187 VSUBS 0.069f
C6737 VOUT.n2188 VSUBS 0.0324f
C6738 VOUT.n2189 VSUBS 0.0365f
C6739 VOUT.n2190 VSUBS 0.0678f
C6740 VOUT.n2191 VSUBS 0.0188f
C6741 VOUT.n2192 VSUBS 0.00925f
C6742 VOUT.n2193 VSUBS 0.0373f
C6743 VOUT.n2194 VSUBS 0.223f
C6744 VOUT.n2195 VSUBS 0.223f
C6745 VOUT.t498 VSUBS 0.0294f
C6746 VOUT.t133 VSUBS 0.0294f
C6747 VOUT.n2196 VSUBS 0.069f
C6748 VOUT.n2197 VSUBS 0.0324f
C6749 VOUT.n2198 VSUBS 0.0365f
C6750 VOUT.n2199 VSUBS 0.0678f
C6751 VOUT.n2200 VSUBS 0.0188f
C6752 VOUT.n2201 VSUBS 0.00925f
C6753 VOUT.n2202 VSUBS 0.0373f
C6754 VOUT.n2203 VSUBS 0.223f
C6755 VOUT.n2204 VSUBS 0.223f
C6756 VOUT.t462 VSUBS 0.0294f
C6757 VOUT.t3 VSUBS 0.0294f
C6758 VOUT.n2205 VSUBS 0.069f
C6759 VOUT.n2206 VSUBS 0.0324f
C6760 VOUT.n2207 VSUBS 0.0365f
C6761 VOUT.n2208 VSUBS 0.0678f
C6762 VOUT.n2209 VSUBS 0.0188f
C6763 VOUT.n2210 VSUBS 0.00925f
C6764 VOUT.n2211 VSUBS 0.0373f
C6765 VOUT.n2212 VSUBS 0.223f
C6766 VOUT.n2213 VSUBS 0.223f
C6767 VOUT.t123 VSUBS 0.0294f
C6768 VOUT.t101 VSUBS 0.0294f
C6769 VOUT.n2214 VSUBS 0.069f
C6770 VOUT.n2215 VSUBS 0.0324f
C6771 VOUT.n2216 VSUBS 0.0365f
C6772 VOUT.n2217 VSUBS 0.0678f
C6773 VOUT.n2218 VSUBS 0.0188f
C6774 VOUT.n2219 VSUBS 0.00925f
C6775 VOUT.n2220 VSUBS 0.0373f
C6776 VOUT.n2221 VSUBS 0.223f
C6777 VOUT.n2222 VSUBS 0.223f
C6778 VOUT.t376 VSUBS 0.0294f
C6779 VOUT.t340 VSUBS 0.0294f
C6780 VOUT.n2223 VSUBS 0.069f
C6781 VOUT.n2224 VSUBS 0.0324f
C6782 VOUT.n2225 VSUBS 0.0365f
C6783 VOUT.n2226 VSUBS 0.0678f
C6784 VOUT.n2227 VSUBS 0.0188f
C6785 VOUT.n2228 VSUBS 0.00925f
C6786 VOUT.n2229 VSUBS 0.0373f
C6787 VOUT.n2230 VSUBS 0.223f
C6788 VOUT.n2231 VSUBS 0.223f
C6789 VOUT.t82 VSUBS 0.0294f
C6790 VOUT.t71 VSUBS 0.0294f
C6791 VOUT.n2232 VSUBS 0.069f
C6792 VOUT.n2233 VSUBS 0.0324f
C6793 VOUT.n2234 VSUBS 0.0365f
C6794 VOUT.n2235 VSUBS 0.0678f
C6795 VOUT.n2236 VSUBS 0.0188f
C6796 VOUT.n2237 VSUBS 0.00925f
C6797 VOUT.n2238 VSUBS 0.0373f
C6798 VOUT.n2239 VSUBS 0.223f
C6799 VOUT.n2240 VSUBS 0.223f
C6800 VOUT.t44 VSUBS 0.0294f
C6801 VOUT.t381 VSUBS 0.0294f
C6802 VOUT.n2241 VSUBS 0.069f
C6803 VOUT.n2242 VSUBS 0.0324f
C6804 VOUT.n2243 VSUBS 0.0365f
C6805 VOUT.n2244 VSUBS 0.0678f
C6806 VOUT.n2245 VSUBS 0.0188f
C6807 VOUT.n2246 VSUBS 0.00925f
C6808 VOUT.n2247 VSUBS 0.0373f
C6809 VOUT.n2248 VSUBS 0.223f
C6810 VOUT.n2249 VSUBS 0.223f
C6811 VOUT.t425 VSUBS 0.0294f
C6812 VOUT.n2250 VSUBS 0.0984f
C6813 VOUT.n2251 VSUBS 0.0324f
C6814 VOUT.n2252 VSUBS 0.0365f
C6815 VOUT.n2253 VSUBS 0.0678f
C6816 VOUT.n2254 VSUBS 0.0188f
C6817 VOUT.n2255 VSUBS 0.00925f
C6818 VOUT.n2256 VSUBS 0.0373f
C6819 VOUT.n2257 VSUBS 0.119f
C6820 VOUT.t8 VSUBS 0.0294f
C6821 VOUT.n2258 VSUBS 0.0985f
C6822 VOUT.n2259 VSUBS 0.0338f
C6823 VOUT.n2260 VSUBS 0.0365f
C6824 VOUT.n2261 VSUBS 0.0707f
C6825 VOUT.n2262 VSUBS 0.0184f
C6826 VOUT.n2263 VSUBS 0.00899f
C6827 VOUT.n2264 VSUBS 0.0373f
C6828 VOUT.t496 VSUBS 0.0294f
C6829 VOUT.t32 VSUBS 0.0294f
C6830 VOUT.n2265 VSUBS 0.0691f
C6831 VOUT.n2266 VSUBS 0.0338f
C6832 VOUT.n2267 VSUBS 0.0365f
C6833 VOUT.n2268 VSUBS 0.0707f
C6834 VOUT.n2269 VSUBS 0.0184f
C6835 VOUT.n2270 VSUBS 0.00899f
C6836 VOUT.n2271 VSUBS 0.0373f
C6837 VOUT.t80 VSUBS 0.0294f
C6838 VOUT.t505 VSUBS 0.0294f
C6839 VOUT.n2272 VSUBS 0.0691f
C6840 VOUT.n2273 VSUBS 0.0338f
C6841 VOUT.n2274 VSUBS 0.0365f
C6842 VOUT.n2275 VSUBS 0.0707f
C6843 VOUT.n2276 VSUBS 0.0184f
C6844 VOUT.n2277 VSUBS 0.00899f
C6845 VOUT.n2278 VSUBS 0.0373f
C6846 VOUT.t507 VSUBS 0.0294f
C6847 VOUT.t363 VSUBS 0.0294f
C6848 VOUT.n2279 VSUBS 0.0691f
C6849 VOUT.n2280 VSUBS 0.0338f
C6850 VOUT.n2281 VSUBS 0.0365f
C6851 VOUT.n2282 VSUBS 0.0707f
C6852 VOUT.n2283 VSUBS 0.0184f
C6853 VOUT.n2284 VSUBS 0.00899f
C6854 VOUT.n2285 VSUBS 0.0373f
C6855 VOUT.t125 VSUBS 0.0294f
C6856 VOUT.t378 VSUBS 0.0294f
C6857 VOUT.n2286 VSUBS 0.0691f
C6858 VOUT.n2287 VSUBS 0.0338f
C6859 VOUT.n2288 VSUBS 0.0365f
C6860 VOUT.n2289 VSUBS 0.0707f
C6861 VOUT.n2290 VSUBS 0.0184f
C6862 VOUT.n2291 VSUBS 0.00899f
C6863 VOUT.n2292 VSUBS 0.0373f
C6864 VOUT.t65 VSUBS 0.0294f
C6865 VOUT.t12 VSUBS 0.0294f
C6866 VOUT.n2293 VSUBS 0.0691f
C6867 VOUT.n2294 VSUBS 0.0338f
C6868 VOUT.n2295 VSUBS 0.0365f
C6869 VOUT.n2296 VSUBS 0.0707f
C6870 VOUT.n2297 VSUBS 0.0184f
C6871 VOUT.n2298 VSUBS 0.00899f
C6872 VOUT.n2299 VSUBS 0.0373f
C6873 VOUT.t20 VSUBS 0.0294f
C6874 VOUT.t112 VSUBS 0.0294f
C6875 VOUT.n2300 VSUBS 0.0691f
C6876 VOUT.n2301 VSUBS 0.0338f
C6877 VOUT.n2302 VSUBS 0.0365f
C6878 VOUT.n2303 VSUBS 0.0707f
C6879 VOUT.n2304 VSUBS 0.0184f
C6880 VOUT.n2305 VSUBS 0.00899f
C6881 VOUT.n2306 VSUBS 0.0373f
C6882 VOUT.t70 VSUBS 0.0294f
C6883 VOUT.t58 VSUBS 0.0294f
C6884 VOUT.n2307 VSUBS 0.0691f
C6885 VOUT.n2308 VSUBS 0.0338f
C6886 VOUT.n2309 VSUBS 0.0365f
C6887 VOUT.n2310 VSUBS 0.0707f
C6888 VOUT.n2311 VSUBS 0.0184f
C6889 VOUT.n2312 VSUBS 0.00899f
C6890 VOUT.n2313 VSUBS 0.0373f
C6891 VOUT.t39 VSUBS 0.0294f
C6892 VOUT.t111 VSUBS 0.0294f
C6893 VOUT.n2314 VSUBS 0.0691f
C6894 VOUT.n2315 VSUBS 0.0338f
C6895 VOUT.n2316 VSUBS 0.0365f
C6896 VOUT.n2317 VSUBS 0.0707f
C6897 VOUT.n2318 VSUBS 0.0184f
C6898 VOUT.n2319 VSUBS 0.00899f
C6899 VOUT.n2320 VSUBS 0.0373f
C6900 VOUT.t352 VSUBS 0.0294f
C6901 VOUT.t509 VSUBS 0.0294f
C6902 VOUT.n2321 VSUBS 0.0691f
C6903 VOUT.n2322 VSUBS 0.0338f
C6904 VOUT.n2323 VSUBS 0.0365f
C6905 VOUT.n2324 VSUBS 0.0707f
C6906 VOUT.n2325 VSUBS 0.0184f
C6907 VOUT.n2326 VSUBS 0.00899f
C6908 VOUT.n2327 VSUBS 0.0373f
C6909 VOUT.t508 VSUBS 0.0294f
C6910 VOUT.t373 VSUBS 0.0294f
C6911 VOUT.n2328 VSUBS 0.0691f
C6912 VOUT.n2329 VSUBS 0.0338f
C6913 VOUT.n2330 VSUBS 0.0365f
C6914 VOUT.n2331 VSUBS 0.0707f
C6915 VOUT.n2332 VSUBS 0.0184f
C6916 VOUT.n2333 VSUBS 0.00899f
C6917 VOUT.n2334 VSUBS 0.0373f
C6918 VOUT.t107 VSUBS 0.0294f
C6919 VOUT.t99 VSUBS 0.0294f
C6920 VOUT.n2335 VSUBS 0.0691f
C6921 VOUT.n2336 VSUBS 0.0338f
C6922 VOUT.n2337 VSUBS 0.0365f
C6923 VOUT.n2338 VSUBS 0.0707f
C6924 VOUT.n2339 VSUBS 0.0184f
C6925 VOUT.n2340 VSUBS 0.00899f
C6926 VOUT.n2341 VSUBS 0.0373f
C6927 VOUT.t364 VSUBS 0.0294f
C6928 VOUT.t77 VSUBS 0.0294f
C6929 VOUT.n2342 VSUBS 0.0691f
C6930 VOUT.n2343 VSUBS 0.0338f
C6931 VOUT.n2344 VSUBS 0.0365f
C6932 VOUT.n2345 VSUBS 0.0707f
C6933 VOUT.n2346 VSUBS 0.0184f
C6934 VOUT.n2347 VSUBS 0.00899f
C6935 VOUT.n2348 VSUBS 0.0373f
C6936 VOUT.t343 VSUBS 0.0294f
C6937 VOUT.t344 VSUBS 0.0294f
C6938 VOUT.n2349 VSUBS 0.0691f
C6939 VOUT.n2350 VSUBS 0.0338f
C6940 VOUT.n2351 VSUBS 0.0365f
C6941 VOUT.n2352 VSUBS 0.0707f
C6942 VOUT.n2353 VSUBS 0.0184f
C6943 VOUT.n2354 VSUBS 0.00899f
C6944 VOUT.n2355 VSUBS 0.0373f
C6945 VOUT.t86 VSUBS 0.0294f
C6946 VOUT.t367 VSUBS 0.0294f
C6947 VOUT.n2356 VSUBS 0.0691f
C6948 VOUT.n2357 VSUBS 0.0338f
C6949 VOUT.n2358 VSUBS 0.0365f
C6950 VOUT.n2359 VSUBS 0.0707f
C6951 VOUT.n2360 VSUBS 0.0184f
C6952 VOUT.n2361 VSUBS 0.00899f
C6953 VOUT.n2362 VSUBS 0.0373f
C6954 VOUT.t495 VSUBS 0.0294f
C6955 VOUT.t18 VSUBS 0.0294f
C6956 VOUT.n2363 VSUBS 0.0691f
C6957 VOUT.n2364 VSUBS 0.0338f
C6958 VOUT.n2365 VSUBS 0.0365f
C6959 VOUT.n2366 VSUBS 0.0707f
C6960 VOUT.n2367 VSUBS 0.0184f
C6961 VOUT.n2368 VSUBS 0.00899f
C6962 VOUT.n2369 VSUBS 0.0373f
C6963 VOUT.t9 VSUBS 0.0294f
C6964 VOUT.t4 VSUBS 0.0294f
C6965 VOUT.n2370 VSUBS 0.0691f
C6966 VOUT.n2371 VSUBS 0.0338f
C6967 VOUT.n2372 VSUBS 0.0365f
C6968 VOUT.n2373 VSUBS 0.0707f
C6969 VOUT.n2374 VSUBS 0.0184f
C6970 VOUT.n2375 VSUBS 0.00899f
C6971 VOUT.n2376 VSUBS 0.0373f
C6972 VOUT.t405 VSUBS 0.0294f
C6973 VOUT.t83 VSUBS 0.0294f
C6974 VOUT.n2377 VSUBS 0.0691f
C6975 VOUT.n2378 VSUBS 0.0338f
C6976 VOUT.n2379 VSUBS 0.0365f
C6977 VOUT.n2380 VSUBS 0.0707f
C6978 VOUT.n2381 VSUBS 0.0184f
C6979 VOUT.n2382 VSUBS 0.00899f
C6980 VOUT.n2383 VSUBS 0.0373f
C6981 VOUT.t115 VSUBS 0.0294f
C6982 VOUT.t504 VSUBS 0.0294f
C6983 VOUT.n2384 VSUBS 0.0691f
C6984 VOUT.n2385 VSUBS 0.0338f
C6985 VOUT.n2386 VSUBS 0.0365f
C6986 VOUT.n2387 VSUBS 0.0707f
C6987 VOUT.n2388 VSUBS 0.0184f
C6988 VOUT.n2389 VSUBS 0.00899f
C6989 VOUT.n2390 VSUBS 0.0373f
C6990 VOUT.t358 VSUBS 0.0294f
C6991 VOUT.t98 VSUBS 0.0294f
C6992 VOUT.n2391 VSUBS 0.0691f
C6993 VOUT.n2392 VSUBS 0.0338f
C6994 VOUT.n2393 VSUBS 0.0365f
C6995 VOUT.n2394 VSUBS 0.0707f
C6996 VOUT.n2395 VSUBS 0.0184f
C6997 VOUT.n2396 VSUBS 0.00899f
C6998 VOUT.n2397 VSUBS 0.0373f
C6999 VOUT.t365 VSUBS 0.0294f
C7000 VOUT.n2398 VSUBS 0.0985f
C7001 VOUT.n2399 VSUBS 0.0338f
C7002 VOUT.n2400 VSUBS 0.041f
C7003 VOUT.n2401 VSUBS 0.0707f
C7004 VOUT.n2402 VSUBS 0.0184f
C7005 VOUT.n2403 VSUBS 0.00899f
C7006 VOUT.n2404 VSUBS 0.0373f
C7007 VOUT.n2405 VSUBS 0.322f
C7008 VOUT.n2406 VSUBS 0.223f
C7009 VOUT.n2407 VSUBS 0.223f
C7010 VOUT.n2408 VSUBS 0.223f
C7011 VOUT.n2409 VSUBS 0.223f
C7012 VOUT.n2410 VSUBS 0.223f
C7013 VOUT.n2411 VSUBS 0.223f
C7014 VOUT.n2412 VSUBS 0.223f
C7015 VOUT.n2413 VSUBS 0.223f
C7016 VOUT.n2414 VSUBS 0.223f
C7017 VOUT.n2415 VSUBS 0.223f
C7018 VOUT.n2416 VSUBS 0.223f
C7019 VOUT.n2417 VSUBS 0.223f
C7020 VOUT.n2418 VSUBS 0.223f
C7021 VOUT.n2419 VSUBS 0.223f
C7022 VOUT.n2420 VSUBS 0.223f
C7023 VOUT.n2421 VSUBS 0.223f
C7024 VOUT.n2422 VSUBS 0.223f
C7025 VOUT.n2423 VSUBS 0.223f
C7026 VOUT.n2424 VSUBS 0.223f
C7027 VOUT.n2425 VSUBS 0.223f
C7028 VOUT.n2426 VSUBS 0.223f
C7029 VOUT.n2427 VSUBS 0.223f
C7030 VOUT.n2428 VSUBS 0.223f
C7031 VOUT.n2429 VSUBS 0.223f
C7032 VOUT.n2430 VSUBS 0.223f
C7033 VOUT.n2431 VSUBS 0.223f
C7034 VOUT.n2432 VSUBS 0.223f
C7035 VOUT.n2433 VSUBS 0.223f
C7036 VOUT.n2434 VSUBS 0.223f
C7037 VOUT.n2435 VSUBS 0.223f
C7038 VOUT.n2436 VSUBS 0.223f
C7039 VOUT.n2437 VSUBS 0.223f
C7040 VOUT.n2438 VSUBS 0.223f
C7041 VOUT.n2439 VSUBS 0.223f
C7042 VOUT.n2440 VSUBS 0.223f
C7043 VOUT.n2441 VSUBS 0.223f
C7044 VOUT.n2442 VSUBS 0.223f
C7045 VOUT.n2443 VSUBS 0.223f
C7046 VOUT.n2444 VSUBS 0.223f
C7047 VOUT.n2445 VSUBS 0.648f
C7048 VOUT.n2446 VSUBS 1.33f
C7049 VOUT.n2447 VSUBS 1.1f
C7050 VOUT.n2448 VSUBS 1.08f
C7051 VOUT.n2449 VSUBS 2.49f
C7052 VOUT.n2450 VSUBS 7.11f
C7053 VOUT.n2451 VSUBS 1.09f
C7054 VOUT.n2452 VSUBS 1.09f
C7055 VOUT.n2453 VSUBS 1.09f
C7056 VOUT.n2454 VSUBS 2.61f
C7057 VOUT.n2455 VSUBS 5.54f
C7058 VDD.n0 VSUBS 0.0155f
C7059 VDD.n1 VSUBS 0.164f
C7060 VDD.n2 VSUBS 0.0155f
C7061 VDD.n3 VSUBS 0.164f
C7062 VDD.n4 VSUBS 0.0155f
C7063 VDD.n5 VSUBS 0.164f
C7064 VDD.n6 VSUBS 0.0155f
C7065 VDD.n7 VSUBS 0.164f
C7066 VDD.n8 VSUBS 0.0155f
C7067 VDD.n9 VSUBS 0.127f
C7068 VDD.n10 VSUBS 0.0155f
C7069 VDD.n11 VSUBS 0.0448f
C7070 VDD.n12 VSUBS 0.0198f
C7071 VDD.n13 VSUBS 0.0448f
C7072 VDD.n14 VSUBS 0.0155f
C7073 VDD.n15 VSUBS 0.0448f
C7074 VDD.n16 VSUBS 0.0198f
C7075 VDD.n17 VSUBS 0.0448f
C7076 VDD.n18 VSUBS 0.0155f
C7077 VDD.n19 VSUBS 0.0448f
C7078 VDD.n20 VSUBS 0.0198f
C7079 VDD.n21 VSUBS 0.0448f
C7080 VDD.n22 VSUBS 0.0155f
C7081 VDD.n23 VSUBS 0.0448f
C7082 VDD.n24 VSUBS 0.0198f
C7083 VDD.n25 VSUBS 0.0448f
C7084 VDD.n26 VSUBS 0.0155f
C7085 VDD.n27 VSUBS 0.0448f
C7086 VDD.n28 VSUBS 0.0198f
C7087 VDD.n29 VSUBS 0.0448f
C7088 VDD.n30 VSUBS 0.0155f
C7089 VDD.n31 VSUBS 0.0448f
C7090 VDD.n32 VSUBS 0.0198f
C7091 VDD.n33 VSUBS 0.0448f
C7092 VDD.n34 VSUBS 0.0155f
C7093 VDD.n35 VSUBS 0.0448f
C7094 VDD.n36 VSUBS 0.0198f
C7095 VDD.n37 VSUBS 0.0448f
C7096 VDD.n38 VSUBS 0.0155f
C7097 VDD.n39 VSUBS 0.0448f
C7098 VDD.n40 VSUBS 0.0198f
C7099 VDD.n41 VSUBS 0.0448f
C7100 VDD.n42 VSUBS 0.0155f
C7101 VDD.n43 VSUBS 0.0448f
C7102 VDD.n44 VSUBS 0.0198f
C7103 VDD.n45 VSUBS 0.0448f
C7104 VDD.n46 VSUBS 0.0155f
C7105 VDD.n47 VSUBS 0.0448f
C7106 VDD.n48 VSUBS 0.0198f
C7107 VDD.n49 VSUBS 0.0448f
C7108 VDD.n50 VSUBS 0.0155f
C7109 VDD.n51 VSUBS 0.0448f
C7110 VDD.n52 VSUBS 0.0198f
C7111 VDD.n53 VSUBS 0.0448f
C7112 VDD.n54 VSUBS 0.0155f
C7113 VDD.n55 VSUBS 0.0448f
C7114 VDD.n56 VSUBS 0.0198f
C7115 VDD.n57 VSUBS 0.0448f
C7116 VDD.n58 VSUBS 0.0155f
C7117 VDD.n59 VSUBS 0.0448f
C7118 VDD.n60 VSUBS 0.0198f
C7119 VDD.n61 VSUBS 0.0448f
C7120 VDD.n62 VSUBS 0.0155f
C7121 VDD.n63 VSUBS 0.0448f
C7122 VDD.n64 VSUBS 0.0198f
C7123 VDD.n65 VSUBS 0.0448f
C7124 VDD.n66 VSUBS 0.0327f
C7125 VDD.n67 VSUBS 0.0448f
C7126 VDD.n68 VSUBS 0.0198f
C7127 VDD.n69 VSUBS 0.0705f
C7128 VDD.n70 VSUBS 0.0198f
C7129 VDD.n71 VSUBS 0.0896f
C7130 VDD.n72 VSUBS 0.0198f
C7131 VDD.n73 VSUBS 0.0896f
C7132 VDD.n74 VSUBS 0.0198f
C7133 VDD.n75 VSUBS 0.0896f
C7134 VDD.n76 VSUBS 0.0842f
C7135 VDD.n77 VSUBS 0.0198f
C7136 VDD.n78 VSUBS 0.0896f
C7137 VDD.n79 VSUBS 0.0842f
C7138 VDD.n80 VSUBS 0.0198f
C7139 VDD.n81 VSUBS 0.0652f
C7140 VDD.n82 VSUBS 0.0842f
C7141 VDD.n83 VSUBS 0.0198f
C7142 VDD.n84 VSUBS 0.0619f
C7143 VDD.n85 VSUBS 0.142f
C7144 VDD.n86 VSUBS 0.0325f
C7145 VDD.n87 VSUBS 0.18f
C7146 VDD.n88 VSUBS 0.0155f
C7147 VDD.n89 VSUBS 0.119f
C7148 VDD.n90 VSUBS 0.358f
C7149 VDD.n91 VSUBS 0.0079f
C7150 VDD.n92 VSUBS 0.0129f
C7151 VDD.n93 VSUBS 0.00241f
C7152 VDD.n94 VSUBS 0.00114f
C7153 VDD.n95 VSUBS 0.00291f
C7154 VDD.n96 VSUBS 6.8e-19
C7155 VDD.n97 VSUBS 0.00393f
C7156 VDD.n98 VSUBS 0.0077f
C7157 VDD.n99 VSUBS 0.00752f
C7158 VDD.n100 VSUBS 0.00376f
C7159 VDD.n101 VSUBS 6.8e-19
C7160 VDD.n102 VSUBS 0.00468f
C7161 VDD.n103 VSUBS 0.00241f
C7162 VDD.n104 VSUBS 0.00114f
C7163 VDD.n105 VSUBS 0.00291f
C7164 VDD.t36 VSUBS 0.0114f
C7165 VDD.n106 VSUBS 0.0345f
C7166 VDD.n107 VSUBS 0.00793f
C7167 VDD.n108 VSUBS 0.013f
C7168 VDD.n109 VSUBS 0.0269f
C7169 VDD.n110 VSUBS 0.00908f
C7170 VDD.n111 VSUBS 0.00929f
C7171 VDD.n112 VSUBS 0.00496f
C7172 VDD.n113 VSUBS 0.00475f
C7173 VDD.n114 VSUBS 0.0828f
C7174 VDD.n115 VSUBS 0.0174f
C7175 VDD.n116 VSUBS 0.0207f
C7176 VDD.n117 VSUBS 0.0842f
C7177 VDD.n118 VSUBS 0.0198f
C7178 VDD.n119 VSUBS 0.0107f
C7179 VDD.n120 VSUBS 0.0114f
C7180 VDD.n121 VSUBS 0.0174f
C7181 VDD.n122 VSUBS 0.032f
C7182 VDD.n124 VSUBS 0.0139f
C7183 VDD.n126 VSUBS 0.0214f
C7184 VDD.n127 VSUBS 0.0174f
C7185 VDD.n128 VSUBS 0.0207f
C7186 VDD.n129 VSUBS 0.0842f
C7187 VDD.n130 VSUBS 0.0198f
C7188 VDD.n131 VSUBS 0.0107f
C7189 VDD.n132 VSUBS 0.0114f
C7190 VDD.n133 VSUBS 0.0174f
C7191 VDD.n134 VSUBS 0.208f
C7192 VDD.n135 VSUBS 0.0384f
C7193 VDD.n136 VSUBS 0.0384f
C7194 VDD.n137 VSUBS 0.0384f
C7195 VDD.n138 VSUBS 0.0277f
C7196 VDD.n139 VSUBS 0.23f
C7197 VDD.n140 VSUBS 0.0321f
C7198 VDD.n141 VSUBS 0.0625f
C7199 VDD.n142 VSUBS 0.0259f
C7200 VDD.n143 VSUBS 0.0388f
C7201 VDD.n144 VSUBS 0.0387f
C7202 VDD.n145 VSUBS 0.0384f
C7203 VDD.t23 VSUBS 0.0095f
C7204 VDD.n146 VSUBS 0.0293f
C7205 VDD.n147 VSUBS 0.0832f
C7206 VDD.n148 VSUBS 0.0438f
C7207 VDD.n149 VSUBS 0.0321f
C7208 VDD.n150 VSUBS 0.0331f
C7209 VDD.n151 VSUBS 0.0321f
C7210 VDD.n152 VSUBS 0.033f
C7211 VDD.n153 VSUBS 0.0232f
C7212 VDD.n154 VSUBS 0.0161f
C7213 VDD.n155 VSUBS 0.0192f
C7214 VDD.n156 VSUBS 0.0298f
C7215 VDD.n157 VSUBS 0.0821f
C7216 VDD.n158 VSUBS 0.351f
C7217 VDD.n159 VSUBS 0.0174f
C7218 VDD.n160 VSUBS 0.0198f
C7219 VDD.n161 VSUBS 0.0398f
C7220 VDD.n162 VSUBS 0.0227f
C7221 VDD.n163 VSUBS 0.0842f
C7222 VDD.n164 VSUBS 0.0198f
C7223 VDD.n165 VSUBS 0.0234f
C7224 VDD.n166 VSUBS 0.0221f
C7225 VDD.n167 VSUBS 0.0842f
C7226 VDD.n168 VSUBS 0.0198f
C7227 VDD.n169 VSUBS 0.0234f
C7228 VDD.n170 VSUBS 0.0842f
C7229 VDD.n171 VSUBS 0.0198f
C7230 VDD.n172 VSUBS 0.0441f
C7231 VDD.n173 VSUBS 0.0842f
C7232 VDD.n174 VSUBS 0.0198f
C7233 VDD.n175 VSUBS 0.0266f
C7234 VDD.n176 VSUBS 0.0229f
C7235 VDD.n177 VSUBS 0.0842f
C7236 VDD.n178 VSUBS 0.0198f
C7237 VDD.n179 VSUBS 0.0234f
C7238 VDD.n180 VSUBS 0.0221f
C7239 VDD.n181 VSUBS 0.0996f
C7240 VDD.n182 VSUBS 0.0842f
C7241 VDD.n183 VSUBS 0.0198f
C7242 VDD.n184 VSUBS 0.0234f
C7243 VDD.n185 VSUBS 0.0221f
C7244 VDD.n186 VSUBS 0.0391f
C7245 VDD.n187 VSUBS 0.0842f
C7246 VDD.n188 VSUBS 0.0198f
C7247 VDD.n189 VSUBS 0.0234f
C7248 VDD.n190 VSUBS 0.0221f
C7249 VDD.n191 VSUBS 0.0391f
C7250 VDD.n192 VSUBS 0.0842f
C7251 VDD.n193 VSUBS 0.0198f
C7252 VDD.n194 VSUBS 0.0234f
C7253 VDD.n195 VSUBS 0.0221f
C7254 VDD.n196 VSUBS 0.0391f
C7255 VDD.n197 VSUBS 0.0842f
C7256 VDD.n198 VSUBS 0.0198f
C7257 VDD.n199 VSUBS 0.0234f
C7258 VDD.n200 VSUBS 0.0842f
C7259 VDD.n201 VSUBS 0.0198f
C7260 VDD.n202 VSUBS 0.0234f
C7261 VDD.n203 VSUBS 0.0221f
C7262 VDD.n204 VSUBS 0.0391f
C7263 VDD.n205 VSUBS 0.0842f
C7264 VDD.n206 VSUBS 0.0198f
C7265 VDD.n207 VSUBS 0.0234f
C7266 VDD.n208 VSUBS 0.0221f
C7267 VDD.n209 VSUBS 0.0391f
C7268 VDD.n210 VSUBS 0.0842f
C7269 VDD.n211 VSUBS 0.0198f
C7270 VDD.n212 VSUBS 0.0234f
C7271 VDD.n213 VSUBS 0.0221f
C7272 VDD.n214 VSUBS 0.0391f
C7273 VDD.n215 VSUBS 0.0842f
C7274 VDD.n216 VSUBS 0.0198f
C7275 VDD.n217 VSUBS 0.0234f
C7276 VDD.n218 VSUBS 0.0221f
C7277 VDD.n219 VSUBS 0.0391f
C7278 VDD.n220 VSUBS 0.0842f
C7279 VDD.n221 VSUBS 0.0198f
C7280 VDD.n222 VSUBS 0.0234f
C7281 VDD.n223 VSUBS 0.0221f
C7282 VDD.n224 VSUBS 0.0391f
C7283 VDD.n225 VSUBS 0.0842f
C7284 VDD.n226 VSUBS 0.0198f
C7285 VDD.n227 VSUBS 0.0234f
C7286 VDD.n228 VSUBS 0.0221f
C7287 VDD.n229 VSUBS 0.0391f
C7288 VDD.n230 VSUBS 0.0842f
C7289 VDD.n231 VSUBS 0.0198f
C7290 VDD.n232 VSUBS 0.0234f
C7291 VDD.n233 VSUBS 0.0221f
C7292 VDD.n234 VSUBS 0.0391f
C7293 VDD.n235 VSUBS 0.0842f
C7294 VDD.n236 VSUBS 0.0198f
C7295 VDD.n237 VSUBS 0.0234f
C7296 VDD.n238 VSUBS 0.0221f
C7297 VDD.n239 VSUBS 0.0391f
C7298 VDD.n240 VSUBS 0.0842f
C7299 VDD.n241 VSUBS 0.0198f
C7300 VDD.n242 VSUBS 0.0227f
C7301 VDD.n243 VSUBS 0.0221f
C7302 VDD.n244 VSUBS 0.0391f
C7303 VDD.n245 VSUBS 0.0842f
C7304 VDD.n246 VSUBS 0.0198f
C7305 VDD.n247 VSUBS 0.0227f
C7306 VDD.n248 VSUBS 0.0221f
C7307 VDD.n249 VSUBS 0.0391f
C7308 VDD.n250 VSUBS 0.0842f
C7309 VDD.n251 VSUBS 0.0198f
C7310 VDD.n252 VSUBS 0.0234f
C7311 VDD.n253 VSUBS 0.0221f
C7312 VDD.n254 VSUBS 0.0391f
C7313 VDD.n255 VSUBS 0.0842f
C7314 VDD.n256 VSUBS 0.0198f
C7315 VDD.n257 VSUBS 0.0234f
C7316 VDD.n258 VSUBS 0.0221f
C7317 VDD.n259 VSUBS 0.0391f
C7318 VDD.n260 VSUBS 0.0985f
C7319 VDD.n261 VSUBS 0.0229f
C7320 VDD.n262 VSUBS 0.0842f
C7321 VDD.n263 VSUBS 0.0198f
C7322 VDD.n264 VSUBS 0.0383f
C7323 VDD.n265 VSUBS 0.0842f
C7324 VDD.n266 VSUBS 0.0198f
C7325 VDD.n267 VSUBS 0.0441f
C7326 VDD.n268 VSUBS 0.0842f
C7327 VDD.n269 VSUBS 0.0198f
C7328 VDD.n270 VSUBS 0.0441f
C7329 VDD.n271 VSUBS 0.0842f
C7330 VDD.n272 VSUBS 0.0198f
C7331 VDD.n273 VSUBS 0.0441f
C7332 VDD.n274 VSUBS 0.0842f
C7333 VDD.n275 VSUBS 0.0198f
C7334 VDD.n276 VSUBS 0.0441f
C7335 VDD.n277 VSUBS 0.0842f
C7336 VDD.n278 VSUBS 0.0198f
C7337 VDD.n279 VSUBS 0.0441f
C7338 VDD.n280 VSUBS 0.0842f
C7339 VDD.n281 VSUBS 0.0198f
C7340 VDD.n282 VSUBS 0.0441f
C7341 VDD.n283 VSUBS 0.0842f
C7342 VDD.n284 VSUBS 0.0198f
C7343 VDD.n285 VSUBS 0.0441f
C7344 VDD.n286 VSUBS 0.0842f
C7345 VDD.n287 VSUBS 0.0198f
C7346 VDD.n288 VSUBS 0.0419f
C7347 VDD.n289 VSUBS 0.0842f
C7348 VDD.n290 VSUBS 0.0198f
C7349 VDD.n291 VSUBS 0.0234f
C7350 VDD.n292 VSUBS 0.023f
C7351 VDD.n293 VSUBS 0.0842f
C7352 VDD.n294 VSUBS 0.0198f
C7353 VDD.n295 VSUBS 0.023f
C7354 VDD.n296 VSUBS 0.0221f
C7355 VDD.n297 VSUBS 0.105f
C7356 VDD.n298 VSUBS 0.0842f
C7357 VDD.n299 VSUBS 0.0198f
C7358 VDD.n300 VSUBS 0.0224f
C7359 VDD.n301 VSUBS 0.0221f
C7360 VDD.n302 VSUBS 0.0391f
C7361 VDD.n303 VSUBS 0.0842f
C7362 VDD.n304 VSUBS 0.0198f
C7363 VDD.n305 VSUBS 0.0234f
C7364 VDD.n306 VSUBS 0.0221f
C7365 VDD.n307 VSUBS 0.0391f
C7366 VDD.n308 VSUBS 0.0842f
C7367 VDD.n309 VSUBS 0.0198f
C7368 VDD.n310 VSUBS 0.0234f
C7369 VDD.n311 VSUBS 0.0221f
C7370 VDD.n312 VSUBS 0.0391f
C7371 VDD.n313 VSUBS 0.0842f
C7372 VDD.n314 VSUBS 0.0198f
C7373 VDD.n315 VSUBS 0.0234f
C7374 VDD.n316 VSUBS 0.0221f
C7375 VDD.n317 VSUBS 0.0391f
C7376 VDD.n318 VSUBS 0.0842f
C7377 VDD.n319 VSUBS 0.0198f
C7378 VDD.n320 VSUBS 0.0234f
C7379 VDD.n321 VSUBS 0.0221f
C7380 VDD.n322 VSUBS 0.0391f
C7381 VDD.n323 VSUBS 0.0842f
C7382 VDD.n324 VSUBS 0.0198f
C7383 VDD.n325 VSUBS 0.0234f
C7384 VDD.n326 VSUBS 0.0221f
C7385 VDD.n327 VSUBS 0.0391f
C7386 VDD.n328 VSUBS 0.0842f
C7387 VDD.n329 VSUBS 0.0198f
C7388 VDD.n330 VSUBS 0.0234f
C7389 VDD.n331 VSUBS 0.0221f
C7390 VDD.n332 VSUBS 0.0391f
C7391 VDD.n333 VSUBS 0.0842f
C7392 VDD.n334 VSUBS 0.0198f
C7393 VDD.n335 VSUBS 0.0234f
C7394 VDD.n336 VSUBS 0.0221f
C7395 VDD.n337 VSUBS 0.0391f
C7396 VDD.n338 VSUBS 0.0842f
C7397 VDD.n339 VSUBS 0.0198f
C7398 VDD.n340 VSUBS 0.0234f
C7399 VDD.n341 VSUBS 0.0842f
C7400 VDD.n342 VSUBS 0.0198f
C7401 VDD.n343 VSUBS 0.0234f
C7402 VDD.n344 VSUBS 0.0221f
C7403 VDD.n345 VSUBS 0.0391f
C7404 VDD.n346 VSUBS 0.0842f
C7405 VDD.n347 VSUBS 0.0198f
C7406 VDD.n348 VSUBS 0.0234f
C7407 VDD.n349 VSUBS 0.0221f
C7408 VDD.n350 VSUBS 0.0391f
C7409 VDD.n351 VSUBS 0.0793f
C7410 VDD.n352 VSUBS 0.0198f
C7411 VDD.n353 VSUBS 0.0234f
C7412 VDD.n354 VSUBS 0.0221f
C7413 VDD.n355 VSUBS 0.0391f
C7414 VDD.n356 VSUBS 0.161f
C7415 VDD.n358 VSUBS 0.0198f
C7416 VDD.n359 VSUBS 0.0295f
C7417 VDD.n360 VSUBS 0.0221f
C7418 VDD.n361 VSUBS 0.0494f
C7419 VDD.n362 VSUBS 0.0198f
C7420 VDD.n363 VSUBS 0.0386f
C7421 VDD.n364 VSUBS 0.0333f
C7422 VDD.n365 VSUBS 0.00713f
C7423 VDD.n366 VSUBS 0.0221f
C7424 VDD.n367 VSUBS 0.0781f
C7425 VDD.n368 VSUBS 0.0849f
C7426 VDD.n369 VSUBS 0.0564f
C7427 VDD.n370 VSUBS 0.0287f
C7428 VDD.n371 VSUBS 0.0842f
C7429 VDD.n372 VSUBS 0.0198f
C7430 VDD.n373 VSUBS 0.00447f
C7431 VDD.n374 VSUBS 0.0535f
C7432 VDD.n375 VSUBS 0.0206f
C7433 VDD.n376 VSUBS 0.0391f
C7434 VDD.n377 VSUBS 0.0842f
C7435 VDD.n378 VSUBS 0.0198f
C7436 VDD.n379 VSUBS 0.0228f
C7437 VDD.n380 VSUBS 0.0215f
C7438 VDD.n381 VSUBS 0.0391f
C7439 VDD.n382 VSUBS 0.0842f
C7440 VDD.n383 VSUBS 0.0198f
C7441 VDD.n384 VSUBS 0.0228f
C7442 VDD.n385 VSUBS 0.0215f
C7443 VDD.n386 VSUBS 0.0391f
C7444 VDD.n387 VSUBS 0.0842f
C7445 VDD.n388 VSUBS 0.0198f
C7446 VDD.n389 VSUBS 0.0228f
C7447 VDD.n390 VSUBS 0.0215f
C7448 VDD.n391 VSUBS 0.0391f
C7449 VDD.n392 VSUBS 0.0842f
C7450 VDD.n393 VSUBS 0.0198f
C7451 VDD.n394 VSUBS 0.0228f
C7452 VDD.n395 VSUBS 0.0842f
C7453 VDD.n396 VSUBS 0.0198f
C7454 VDD.n397 VSUBS 0.0228f
C7455 VDD.n398 VSUBS 0.0215f
C7456 VDD.n399 VSUBS 0.0391f
C7457 VDD.n400 VSUBS 0.0842f
C7458 VDD.n401 VSUBS 0.0198f
C7459 VDD.n402 VSUBS 0.0228f
C7460 VDD.n403 VSUBS 0.0215f
C7461 VDD.n404 VSUBS 0.0391f
C7462 VDD.n405 VSUBS 0.0842f
C7463 VDD.n406 VSUBS 0.0198f
C7464 VDD.n407 VSUBS 0.0228f
C7465 VDD.n408 VSUBS 0.0215f
C7466 VDD.n409 VSUBS 0.0391f
C7467 VDD.n410 VSUBS 0.0842f
C7468 VDD.n411 VSUBS 0.0198f
C7469 VDD.n412 VSUBS 0.0228f
C7470 VDD.n413 VSUBS 0.0215f
C7471 VDD.n414 VSUBS 0.0391f
C7472 VDD.n415 VSUBS 0.0842f
C7473 VDD.n416 VSUBS 0.0198f
C7474 VDD.n417 VSUBS 0.0228f
C7475 VDD.n418 VSUBS 0.0215f
C7476 VDD.n419 VSUBS 0.0391f
C7477 VDD.n420 VSUBS 0.0842f
C7478 VDD.n421 VSUBS 0.0198f
C7479 VDD.n422 VSUBS 0.0228f
C7480 VDD.n423 VSUBS 0.0215f
C7481 VDD.n424 VSUBS 0.0391f
C7482 VDD.n425 VSUBS 0.0842f
C7483 VDD.n426 VSUBS 0.0198f
C7484 VDD.n427 VSUBS 0.0228f
C7485 VDD.n428 VSUBS 0.0215f
C7486 VDD.n429 VSUBS 0.0391f
C7487 VDD.n430 VSUBS 0.0842f
C7488 VDD.n431 VSUBS 0.0198f
C7489 VDD.n432 VSUBS 0.0228f
C7490 VDD.n433 VSUBS 0.0215f
C7491 VDD.n434 VSUBS 0.0391f
C7492 VDD.n435 VSUBS 0.0842f
C7493 VDD.n436 VSUBS 0.0198f
C7494 VDD.n437 VSUBS 0.0225f
C7495 VDD.n438 VSUBS 0.0215f
C7496 VDD.n439 VSUBS 0.0391f
C7497 VDD.n440 VSUBS 0.0842f
C7498 VDD.n441 VSUBS 0.0198f
C7499 VDD.n442 VSUBS 0.0218f
C7500 VDD.n443 VSUBS 0.0215f
C7501 VDD.n444 VSUBS 0.0391f
C7502 VDD.n445 VSUBS 0.0842f
C7503 VDD.n446 VSUBS 0.0198f
C7504 VDD.n447 VSUBS 0.0228f
C7505 VDD.n448 VSUBS 0.0215f
C7506 VDD.n449 VSUBS 0.0391f
C7507 VDD.n450 VSUBS 0.0842f
C7508 VDD.n451 VSUBS 0.0198f
C7509 VDD.n452 VSUBS 0.0228f
C7510 VDD.n453 VSUBS 0.0215f
C7511 VDD.n454 VSUBS 0.0391f
C7512 VDD.n455 VSUBS 0.0842f
C7513 VDD.n456 VSUBS 0.0198f
C7514 VDD.n457 VSUBS 0.0228f
C7515 VDD.n458 VSUBS 0.0215f
C7516 VDD.n459 VSUBS 0.0391f
C7517 VDD.n460 VSUBS 0.0842f
C7518 VDD.n461 VSUBS 0.0198f
C7519 VDD.n462 VSUBS 0.0228f
C7520 VDD.n463 VSUBS 0.0215f
C7521 VDD.n464 VSUBS 0.0391f
C7522 VDD.n465 VSUBS 0.0842f
C7523 VDD.n466 VSUBS 0.0198f
C7524 VDD.n467 VSUBS 0.0228f
C7525 VDD.n468 VSUBS 0.0215f
C7526 VDD.n469 VSUBS 0.0391f
C7527 VDD.n470 VSUBS 0.0842f
C7528 VDD.n471 VSUBS 0.0198f
C7529 VDD.n472 VSUBS 0.0228f
C7530 VDD.n473 VSUBS 0.0215f
C7531 VDD.n474 VSUBS 0.0391f
C7532 VDD.n475 VSUBS 0.0842f
C7533 VDD.n476 VSUBS 0.0198f
C7534 VDD.n477 VSUBS 0.0228f
C7535 VDD.n478 VSUBS 0.0215f
C7536 VDD.n479 VSUBS 0.0391f
C7537 VDD.n480 VSUBS 0.0842f
C7538 VDD.n481 VSUBS 0.0198f
C7539 VDD.n482 VSUBS 0.0228f
C7540 VDD.n483 VSUBS 0.0842f
C7541 VDD.n484 VSUBS 0.0198f
C7542 VDD.n485 VSUBS 0.0228f
C7543 VDD.n486 VSUBS 0.0215f
C7544 VDD.n487 VSUBS 0.0391f
C7545 VDD.n488 VSUBS 0.0842f
C7546 VDD.n489 VSUBS 0.0198f
C7547 VDD.n490 VSUBS 0.0228f
C7548 VDD.n491 VSUBS 0.0215f
C7549 VDD.n492 VSUBS 0.0391f
C7550 VDD.n493 VSUBS 0.0842f
C7551 VDD.n494 VSUBS 0.0198f
C7552 VDD.n495 VSUBS 0.0228f
C7553 VDD.n496 VSUBS 0.0215f
C7554 VDD.n497 VSUBS 0.0391f
C7555 VDD.n498 VSUBS 0.0842f
C7556 VDD.n499 VSUBS 0.0198f
C7557 VDD.n500 VSUBS 0.0228f
C7558 VDD.n501 VSUBS 0.0215f
C7559 VDD.n502 VSUBS 0.0391f
C7560 VDD.n503 VSUBS 0.0842f
C7561 VDD.n504 VSUBS 0.0198f
C7562 VDD.n505 VSUBS 0.0228f
C7563 VDD.n506 VSUBS 0.0215f
C7564 VDD.n507 VSUBS 0.0391f
C7565 VDD.n508 VSUBS 0.0842f
C7566 VDD.n509 VSUBS 0.0198f
C7567 VDD.n510 VSUBS 0.0228f
C7568 VDD.n511 VSUBS 0.0215f
C7569 VDD.n512 VSUBS 0.0391f
C7570 VDD.n513 VSUBS 0.0842f
C7571 VDD.n514 VSUBS 0.0198f
C7572 VDD.n515 VSUBS 0.0228f
C7573 VDD.n516 VSUBS 0.0215f
C7574 VDD.n517 VSUBS 0.0391f
C7575 VDD.n518 VSUBS 0.0842f
C7576 VDD.n519 VSUBS 0.0198f
C7577 VDD.n520 VSUBS 0.0228f
C7578 VDD.n521 VSUBS 0.0215f
C7579 VDD.n522 VSUBS 0.0391f
C7580 VDD.n523 VSUBS 0.0842f
C7581 VDD.n524 VSUBS 0.0198f
C7582 VDD.n525 VSUBS 0.0225f
C7583 VDD.n526 VSUBS 0.0215f
C7584 VDD.n527 VSUBS 0.0391f
C7585 VDD.n528 VSUBS 0.0842f
C7586 VDD.n529 VSUBS 0.0198f
C7587 VDD.n530 VSUBS 0.0218f
C7588 VDD.n531 VSUBS 0.0215f
C7589 VDD.n532 VSUBS 0.0391f
C7590 VDD.n533 VSUBS 0.0842f
C7591 VDD.n534 VSUBS 0.0198f
C7592 VDD.n535 VSUBS 0.0228f
C7593 VDD.n536 VSUBS 0.0215f
C7594 VDD.n537 VSUBS 0.0391f
C7595 VDD.n538 VSUBS 0.0842f
C7596 VDD.n539 VSUBS 0.0198f
C7597 VDD.n540 VSUBS 0.0228f
C7598 VDD.n541 VSUBS 0.0215f
C7599 VDD.n542 VSUBS 0.0391f
C7600 VDD.n543 VSUBS 0.0842f
C7601 VDD.n544 VSUBS 0.0198f
C7602 VDD.n545 VSUBS 0.0228f
C7603 VDD.n546 VSUBS 0.0215f
C7604 VDD.n547 VSUBS 0.0391f
C7605 VDD.n548 VSUBS 0.0842f
C7606 VDD.n549 VSUBS 0.0198f
C7607 VDD.n550 VSUBS 0.0228f
C7608 VDD.n551 VSUBS 0.0215f
C7609 VDD.n552 VSUBS 0.0391f
C7610 VDD.n553 VSUBS 0.0842f
C7611 VDD.n554 VSUBS 0.0198f
C7612 VDD.n555 VSUBS 0.0228f
C7613 VDD.n556 VSUBS 0.0215f
C7614 VDD.n557 VSUBS 0.0391f
C7615 VDD.n558 VSUBS 0.0842f
C7616 VDD.n559 VSUBS 0.0198f
C7617 VDD.n560 VSUBS 0.0228f
C7618 VDD.n561 VSUBS 0.0215f
C7619 VDD.n562 VSUBS 0.0391f
C7620 VDD.n563 VSUBS 0.0842f
C7621 VDD.n564 VSUBS 0.0198f
C7622 VDD.n565 VSUBS 0.0228f
C7623 VDD.n566 VSUBS 0.0215f
C7624 VDD.n567 VSUBS 0.0391f
C7625 VDD.n568 VSUBS 0.0842f
C7626 VDD.n569 VSUBS 0.0198f
C7627 VDD.n570 VSUBS 0.0228f
C7628 VDD.n571 VSUBS 0.0842f
C7629 VDD.n572 VSUBS 0.0198f
C7630 VDD.n573 VSUBS 0.0228f
C7631 VDD.n574 VSUBS 0.0215f
C7632 VDD.n575 VSUBS 0.0391f
C7633 VDD.n576 VSUBS 0.0842f
C7634 VDD.n577 VSUBS 0.0198f
C7635 VDD.n578 VSUBS 0.0228f
C7636 VDD.n579 VSUBS 0.0215f
C7637 VDD.n580 VSUBS 0.0391f
C7638 VDD.n581 VSUBS 0.0842f
C7639 VDD.n582 VSUBS 0.0198f
C7640 VDD.n583 VSUBS 0.0228f
C7641 VDD.n584 VSUBS 0.0215f
C7642 VDD.n585 VSUBS 0.0391f
C7643 VDD.n586 VSUBS 0.0842f
C7644 VDD.n587 VSUBS 0.0198f
C7645 VDD.n588 VSUBS 0.0228f
C7646 VDD.n589 VSUBS 0.0215f
C7647 VDD.n590 VSUBS 0.0391f
C7648 VDD.n591 VSUBS 0.0842f
C7649 VDD.n592 VSUBS 0.0198f
C7650 VDD.n593 VSUBS 0.0228f
C7651 VDD.n594 VSUBS 0.0215f
C7652 VDD.n595 VSUBS 0.0391f
C7653 VDD.n596 VSUBS 0.0842f
C7654 VDD.n597 VSUBS 0.0198f
C7655 VDD.n598 VSUBS 0.0228f
C7656 VDD.n599 VSUBS 0.0215f
C7657 VDD.n600 VSUBS 0.0391f
C7658 VDD.n601 VSUBS 0.0842f
C7659 VDD.n602 VSUBS 0.0198f
C7660 VDD.n603 VSUBS 0.0228f
C7661 VDD.n604 VSUBS 0.0215f
C7662 VDD.n605 VSUBS 0.0391f
C7663 VDD.n606 VSUBS 0.0842f
C7664 VDD.n607 VSUBS 0.0198f
C7665 VDD.n608 VSUBS 0.0228f
C7666 VDD.n609 VSUBS 0.0215f
C7667 VDD.n610 VSUBS 0.0391f
C7668 VDD.n611 VSUBS 0.0842f
C7669 VDD.n612 VSUBS 0.0198f
C7670 VDD.n613 VSUBS 0.0225f
C7671 VDD.n614 VSUBS 0.0215f
C7672 VDD.n615 VSUBS 0.0391f
C7673 VDD.n616 VSUBS 0.0842f
C7674 VDD.n617 VSUBS 0.0198f
C7675 VDD.n618 VSUBS 0.0218f
C7676 VDD.n619 VSUBS 0.0215f
C7677 VDD.n620 VSUBS 0.0391f
C7678 VDD.n621 VSUBS 0.0842f
C7679 VDD.n622 VSUBS 0.0198f
C7680 VDD.n623 VSUBS 0.0228f
C7681 VDD.n624 VSUBS 0.0215f
C7682 VDD.n625 VSUBS 0.0391f
C7683 VDD.n626 VSUBS 0.0842f
C7684 VDD.n627 VSUBS 0.0198f
C7685 VDD.n628 VSUBS 0.0228f
C7686 VDD.n629 VSUBS 0.0215f
C7687 VDD.n630 VSUBS 0.0391f
C7688 VDD.n631 VSUBS 0.0842f
C7689 VDD.n632 VSUBS 0.0198f
C7690 VDD.n633 VSUBS 0.0228f
C7691 VDD.n634 VSUBS 0.0215f
C7692 VDD.n635 VSUBS 0.0391f
C7693 VDD.n636 VSUBS 0.0842f
C7694 VDD.n637 VSUBS 0.0198f
C7695 VDD.n638 VSUBS 0.0228f
C7696 VDD.n639 VSUBS 0.0215f
C7697 VDD.n640 VSUBS 0.0391f
C7698 VDD.n641 VSUBS 0.0842f
C7699 VDD.n642 VSUBS 0.0198f
C7700 VDD.n643 VSUBS 0.0228f
C7701 VDD.n644 VSUBS 0.0215f
C7702 VDD.n645 VSUBS 0.0391f
C7703 VDD.n646 VSUBS 0.0842f
C7704 VDD.n647 VSUBS 0.0198f
C7705 VDD.n648 VSUBS 0.0228f
C7706 VDD.n649 VSUBS 0.0215f
C7707 VDD.n650 VSUBS 0.0391f
C7708 VDD.n651 VSUBS 0.0842f
C7709 VDD.n652 VSUBS 0.0198f
C7710 VDD.n653 VSUBS 0.0228f
C7711 VDD.n654 VSUBS 0.0215f
C7712 VDD.n655 VSUBS 0.0391f
C7713 VDD.n656 VSUBS 0.0842f
C7714 VDD.n657 VSUBS 0.0198f
C7715 VDD.n658 VSUBS 0.0228f
C7716 VDD.n659 VSUBS 0.0842f
C7717 VDD.n660 VSUBS 0.0198f
C7718 VDD.n661 VSUBS 0.0228f
C7719 VDD.n662 VSUBS 0.0215f
C7720 VDD.n663 VSUBS 0.0391f
C7721 VDD.n664 VSUBS 0.0842f
C7722 VDD.n665 VSUBS 0.0198f
C7723 VDD.n666 VSUBS 0.0228f
C7724 VDD.n667 VSUBS 0.0215f
C7725 VDD.n668 VSUBS 0.0391f
C7726 VDD.n669 VSUBS 0.0842f
C7727 VDD.n670 VSUBS 0.0198f
C7728 VDD.n671 VSUBS 0.0228f
C7729 VDD.n672 VSUBS 0.0215f
C7730 VDD.n673 VSUBS 0.0391f
C7731 VDD.n674 VSUBS 0.0842f
C7732 VDD.n675 VSUBS 0.0198f
C7733 VDD.n676 VSUBS 0.0228f
C7734 VDD.n677 VSUBS 0.0215f
C7735 VDD.n678 VSUBS 0.0391f
C7736 VDD.n679 VSUBS 0.0842f
C7737 VDD.n680 VSUBS 0.0198f
C7738 VDD.n681 VSUBS 0.0228f
C7739 VDD.n682 VSUBS 0.0215f
C7740 VDD.n683 VSUBS 0.0391f
C7741 VDD.n684 VSUBS 0.0842f
C7742 VDD.n685 VSUBS 0.0198f
C7743 VDD.n686 VSUBS 0.0228f
C7744 VDD.n687 VSUBS 0.0215f
C7745 VDD.n688 VSUBS 0.0391f
C7746 VDD.n689 VSUBS 0.0842f
C7747 VDD.n690 VSUBS 0.0198f
C7748 VDD.n691 VSUBS 0.0228f
C7749 VDD.n692 VSUBS 0.0215f
C7750 VDD.n693 VSUBS 0.0391f
C7751 VDD.n694 VSUBS 0.0842f
C7752 VDD.n695 VSUBS 0.0198f
C7753 VDD.n696 VSUBS 0.0228f
C7754 VDD.n697 VSUBS 0.0215f
C7755 VDD.n698 VSUBS 0.0391f
C7756 VDD.n699 VSUBS 0.0842f
C7757 VDD.n700 VSUBS 0.0198f
C7758 VDD.n701 VSUBS 0.0225f
C7759 VDD.n702 VSUBS 0.0215f
C7760 VDD.n703 VSUBS 0.0391f
C7761 VDD.n704 VSUBS 0.0842f
C7762 VDD.n705 VSUBS 0.0198f
C7763 VDD.n706 VSUBS 0.0218f
C7764 VDD.n707 VSUBS 0.0215f
C7765 VDD.n708 VSUBS 0.0391f
C7766 VDD.n709 VSUBS 0.0842f
C7767 VDD.n710 VSUBS 0.0198f
C7768 VDD.n711 VSUBS 0.0228f
C7769 VDD.n712 VSUBS 0.0215f
C7770 VDD.n713 VSUBS 0.0391f
C7771 VDD.n714 VSUBS 0.0842f
C7772 VDD.n715 VSUBS 0.0198f
C7773 VDD.n716 VSUBS 0.0228f
C7774 VDD.n717 VSUBS 0.0215f
C7775 VDD.n718 VSUBS 0.0391f
C7776 VDD.n719 VSUBS 0.0842f
C7777 VDD.n720 VSUBS 0.0198f
C7778 VDD.n721 VSUBS 0.0228f
C7779 VDD.n722 VSUBS 0.0215f
C7780 VDD.n723 VSUBS 0.0391f
C7781 VDD.n724 VSUBS 0.0842f
C7782 VDD.n725 VSUBS 0.0198f
C7783 VDD.n726 VSUBS 0.0228f
C7784 VDD.n727 VSUBS 0.0215f
C7785 VDD.n728 VSUBS 0.0391f
C7786 VDD.n729 VSUBS 0.0842f
C7787 VDD.n730 VSUBS 0.0198f
C7788 VDD.n731 VSUBS 0.0228f
C7789 VDD.n732 VSUBS 0.0215f
C7790 VDD.n733 VSUBS 0.0391f
C7791 VDD.n734 VSUBS 0.0842f
C7792 VDD.n735 VSUBS 0.0198f
C7793 VDD.n736 VSUBS 0.0228f
C7794 VDD.n737 VSUBS 0.0215f
C7795 VDD.n738 VSUBS 0.0391f
C7796 VDD.n739 VSUBS 0.0842f
C7797 VDD.n740 VSUBS 0.0198f
C7798 VDD.n741 VSUBS 0.0228f
C7799 VDD.n742 VSUBS 0.0215f
C7800 VDD.n743 VSUBS 0.0391f
C7801 VDD.n744 VSUBS 0.0842f
C7802 VDD.n745 VSUBS 0.0198f
C7803 VDD.n746 VSUBS 0.0228f
C7804 VDD.n747 VSUBS 0.0842f
C7805 VDD.n748 VSUBS 0.0198f
C7806 VDD.n749 VSUBS 0.0228f
C7807 VDD.n750 VSUBS 0.0215f
C7808 VDD.n751 VSUBS 0.0391f
C7809 VDD.n752 VSUBS 0.0842f
C7810 VDD.n753 VSUBS 0.0198f
C7811 VDD.n754 VSUBS 0.0228f
C7812 VDD.n755 VSUBS 0.0215f
C7813 VDD.n756 VSUBS 0.0391f
C7814 VDD.n757 VSUBS 0.0842f
C7815 VDD.n758 VSUBS 0.0198f
C7816 VDD.n759 VSUBS 0.0228f
C7817 VDD.n760 VSUBS 0.0215f
C7818 VDD.n761 VSUBS 0.0391f
C7819 VDD.n762 VSUBS 0.0842f
C7820 VDD.n763 VSUBS 0.0198f
C7821 VDD.n764 VSUBS 0.0228f
C7822 VDD.n765 VSUBS 0.0215f
C7823 VDD.n766 VSUBS 0.0391f
C7824 VDD.n767 VSUBS 0.0842f
C7825 VDD.n768 VSUBS 0.0198f
C7826 VDD.n769 VSUBS 0.0228f
C7827 VDD.n770 VSUBS 0.0215f
C7828 VDD.n771 VSUBS 0.0391f
C7829 VDD.n772 VSUBS 0.0842f
C7830 VDD.n773 VSUBS 0.0198f
C7831 VDD.n774 VSUBS 0.0228f
C7832 VDD.n775 VSUBS 0.0215f
C7833 VDD.n776 VSUBS 0.0391f
C7834 VDD.n777 VSUBS 0.0842f
C7835 VDD.n778 VSUBS 0.0198f
C7836 VDD.n779 VSUBS 0.0228f
C7837 VDD.n780 VSUBS 0.0215f
C7838 VDD.n781 VSUBS 0.0391f
C7839 VDD.n782 VSUBS 0.0842f
C7840 VDD.n783 VSUBS 0.0198f
C7841 VDD.n784 VSUBS 0.0228f
C7842 VDD.n785 VSUBS 0.0215f
C7843 VDD.n786 VSUBS 0.0391f
C7844 VDD.n787 VSUBS 0.0842f
C7845 VDD.n788 VSUBS 0.0198f
C7846 VDD.n789 VSUBS 0.0225f
C7847 VDD.n790 VSUBS 0.0215f
C7848 VDD.n791 VSUBS 0.0391f
C7849 VDD.n792 VSUBS 0.0842f
C7850 VDD.n793 VSUBS 0.0198f
C7851 VDD.n794 VSUBS 0.0218f
C7852 VDD.n795 VSUBS 0.0215f
C7853 VDD.n796 VSUBS 0.0391f
C7854 VDD.n797 VSUBS 0.0842f
C7855 VDD.n798 VSUBS 0.0198f
C7856 VDD.n799 VSUBS 0.0228f
C7857 VDD.n800 VSUBS 0.0215f
C7858 VDD.n801 VSUBS 0.0391f
C7859 VDD.n802 VSUBS 0.0842f
C7860 VDD.n803 VSUBS 0.0198f
C7861 VDD.n804 VSUBS 0.0228f
C7862 VDD.n805 VSUBS 0.0215f
C7863 VDD.n806 VSUBS 0.0391f
C7864 VDD.n807 VSUBS 0.0842f
C7865 VDD.n808 VSUBS 0.0198f
C7866 VDD.n809 VSUBS 0.0228f
C7867 VDD.n810 VSUBS 0.0215f
C7868 VDD.n811 VSUBS 0.0391f
C7869 VDD.n812 VSUBS 0.0842f
C7870 VDD.n813 VSUBS 0.0198f
C7871 VDD.n814 VSUBS 0.0228f
C7872 VDD.n815 VSUBS 0.0215f
C7873 VDD.n816 VSUBS 0.0391f
C7874 VDD.n817 VSUBS 0.0842f
C7875 VDD.n818 VSUBS 0.0198f
C7876 VDD.n819 VSUBS 0.0228f
C7877 VDD.n820 VSUBS 0.0215f
C7878 VDD.n821 VSUBS 0.0391f
C7879 VDD.n822 VSUBS 0.0842f
C7880 VDD.n823 VSUBS 0.0198f
C7881 VDD.n824 VSUBS 0.0228f
C7882 VDD.n825 VSUBS 0.0215f
C7883 VDD.n826 VSUBS 0.0391f
C7884 VDD.n827 VSUBS 0.0842f
C7885 VDD.n828 VSUBS 0.0198f
C7886 VDD.n829 VSUBS 0.0228f
C7887 VDD.n830 VSUBS 0.0215f
C7888 VDD.n831 VSUBS 0.0391f
C7889 VDD.n832 VSUBS 0.0842f
C7890 VDD.n833 VSUBS 0.0198f
C7891 VDD.n834 VSUBS 0.0228f
C7892 VDD.n835 VSUBS 0.0842f
C7893 VDD.n836 VSUBS 0.0198f
C7894 VDD.n837 VSUBS 0.0228f
C7895 VDD.n838 VSUBS 0.0215f
C7896 VDD.n839 VSUBS 0.0391f
C7897 VDD.n840 VSUBS 0.0842f
C7898 VDD.n841 VSUBS 0.0198f
C7899 VDD.n842 VSUBS 0.0228f
C7900 VDD.n843 VSUBS 0.0215f
C7901 VDD.n844 VSUBS 0.0391f
C7902 VDD.n845 VSUBS 0.0842f
C7903 VDD.n846 VSUBS 0.0198f
C7904 VDD.n847 VSUBS 0.0228f
C7905 VDD.n848 VSUBS 0.0215f
C7906 VDD.n849 VSUBS 0.0391f
C7907 VDD.n850 VSUBS 0.0842f
C7908 VDD.n851 VSUBS 0.0198f
C7909 VDD.n852 VSUBS 0.0228f
C7910 VDD.n853 VSUBS 0.0215f
C7911 VDD.n854 VSUBS 0.0391f
C7912 VDD.n855 VSUBS 0.0842f
C7913 VDD.n856 VSUBS 0.0198f
C7914 VDD.n857 VSUBS 0.0228f
C7915 VDD.n858 VSUBS 0.0215f
C7916 VDD.n859 VSUBS 0.0391f
C7917 VDD.n860 VSUBS 0.0842f
C7918 VDD.n861 VSUBS 0.0198f
C7919 VDD.n862 VSUBS 0.0228f
C7920 VDD.n863 VSUBS 0.0215f
C7921 VDD.n864 VSUBS 0.0391f
C7922 VDD.n865 VSUBS 0.162f
C7923 VDD.n867 VSUBS 0.0333f
C7924 VDD.n868 VSUBS 0.00735f
C7925 VDD.n869 VSUBS 0.0842f
C7926 VDD.n870 VSUBS 0.0198f
C7927 VDD.n871 VSUBS 0.0849f
C7928 VDD.n872 VSUBS 0.0557f
C7929 VDD.n873 VSUBS 0.0287f
C7930 VDD.n874 VSUBS 0.00449f
C7931 VDD.n875 VSUBS 0.0516f
C7932 VDD.n876 VSUBS 0.019f
C7933 VDD.n877 VSUBS 0.0391f
C7934 VDD.n878 VSUBS 0.104f
C7935 VDD.n879 VSUBS 0.0548f
C7936 VDD.n881 VSUBS 0.0198f
C7937 VDD.n882 VSUBS 0.0455f
C7938 VDD.n883 VSUBS 0.0793f
C7939 VDD.n884 VSUBS 0.0198f
C7940 VDD.n885 VSUBS 0.0381f
C7941 VDD.n886 VSUBS 0.0227f
C7942 VDD.n887 VSUBS 0.0842f
C7943 VDD.n888 VSUBS 0.0198f
C7944 VDD.n889 VSUBS 0.00936f
C7945 VDD.n890 VSUBS 0.0127f
C7946 VDD.n891 VSUBS 0.0163f
C7947 VDD.n892 VSUBS 0.327f
C7948 VDD.n893 VSUBS 0.0842f
C7949 VDD.n894 VSUBS 0.0198f
C7950 VDD.n895 VSUBS 0.0227f
C7951 VDD.n896 VSUBS 0.0227f
C7952 VDD.n897 VSUBS 0.0842f
C7953 VDD.n898 VSUBS 0.0198f
C7954 VDD.n899 VSUBS 0.00903f
C7955 VDD.n900 VSUBS 0.0127f
C7956 VDD.n901 VSUBS 0.016f
C7957 VDD.n902 VSUBS 0.0258f
C7958 VDD.n903 VSUBS 0.0227f
C7959 VDD.n904 VSUBS 0.038f
C7960 VDD.n905 VSUBS 0.0842f
C7961 VDD.n906 VSUBS 0.0198f
C7962 VDD.n907 VSUBS 0.0241f
C7963 VDD.n908 VSUBS 0.0227f
C7964 VDD.n909 VSUBS 0.0391f
C7965 VDD.n910 VSUBS 0.0842f
C7966 VDD.n911 VSUBS 0.0198f
C7967 VDD.n912 VSUBS 0.0241f
C7968 VDD.n913 VSUBS 0.0227f
C7969 VDD.n914 VSUBS 0.0391f
C7970 VDD.n915 VSUBS 0.0842f
C7971 VDD.n916 VSUBS 0.0198f
C7972 VDD.n917 VSUBS 0.0241f
C7973 VDD.n918 VSUBS 0.0842f
C7974 VDD.n919 VSUBS 0.0198f
C7975 VDD.n920 VSUBS 0.0241f
C7976 VDD.n921 VSUBS 0.0227f
C7977 VDD.n922 VSUBS 0.0391f
C7978 VDD.n923 VSUBS 0.0842f
C7979 VDD.n924 VSUBS 0.0198f
C7980 VDD.n925 VSUBS 0.0241f
C7981 VDD.n926 VSUBS 0.0227f
C7982 VDD.n927 VSUBS 0.0391f
C7983 VDD.n928 VSUBS 0.0842f
C7984 VDD.n929 VSUBS 0.0198f
C7985 VDD.n930 VSUBS 0.0241f
C7986 VDD.n931 VSUBS 0.0227f
C7987 VDD.n932 VSUBS 0.0391f
C7988 VDD.n933 VSUBS 0.0842f
C7989 VDD.n934 VSUBS 0.0198f
C7990 VDD.n935 VSUBS 0.0241f
C7991 VDD.n936 VSUBS 0.0227f
C7992 VDD.n937 VSUBS 0.0391f
C7993 VDD.n938 VSUBS 0.0842f
C7994 VDD.n939 VSUBS 0.0198f
C7995 VDD.n940 VSUBS 0.0241f
C7996 VDD.n941 VSUBS 0.0227f
C7997 VDD.n942 VSUBS 0.0391f
C7998 VDD.n943 VSUBS 0.0842f
C7999 VDD.n944 VSUBS 0.0198f
C8000 VDD.n945 VSUBS 0.0241f
C8001 VDD.n946 VSUBS 0.0227f
C8002 VDD.n947 VSUBS 0.0391f
C8003 VDD.n948 VSUBS 0.0842f
C8004 VDD.n949 VSUBS 0.0198f
C8005 VDD.n950 VSUBS 0.0455f
C8006 VDD.n951 VSUBS 0.0842f
C8007 VDD.n952 VSUBS 0.0198f
C8008 VDD.n953 VSUBS 0.0455f
C8009 VDD.n954 VSUBS 0.0842f
C8010 VDD.n955 VSUBS 0.0198f
C8011 VDD.n956 VSUBS 0.0455f
C8012 VDD.n957 VSUBS 0.0842f
C8013 VDD.n958 VSUBS 0.0198f
C8014 VDD.n959 VSUBS 0.0455f
C8015 VDD.n960 VSUBS 0.0842f
C8016 VDD.n961 VSUBS 0.0198f
C8017 VDD.n962 VSUBS 0.0455f
C8018 VDD.n963 VSUBS 0.0842f
C8019 VDD.n964 VSUBS 0.0198f
C8020 VDD.n965 VSUBS 0.0455f
C8021 VDD.n966 VSUBS 0.0842f
C8022 VDD.n967 VSUBS 0.0198f
C8023 VDD.n968 VSUBS 0.0455f
C8024 VDD.n969 VSUBS 0.0842f
C8025 VDD.n970 VSUBS 0.0198f
C8026 VDD.n971 VSUBS 0.0455f
C8027 VDD.n972 VSUBS 0.0842f
C8028 VDD.n973 VSUBS 0.0198f
C8029 VDD.n974 VSUBS 0.0455f
C8030 VDD.n975 VSUBS 0.0842f
C8031 VDD.n976 VSUBS 0.0198f
C8032 VDD.n977 VSUBS 0.0455f
C8033 VDD.n978 VSUBS 0.0842f
C8034 VDD.n979 VSUBS 0.0198f
C8035 VDD.n980 VSUBS 0.0455f
C8036 VDD.n981 VSUBS 0.0842f
C8037 VDD.n982 VSUBS 0.0198f
C8038 VDD.n983 VSUBS 0.0455f
C8039 VDD.n984 VSUBS 0.0842f
C8040 VDD.n985 VSUBS 0.0198f
C8041 VDD.n986 VSUBS 0.0455f
C8042 VDD.n987 VSUBS 0.0842f
C8043 VDD.n988 VSUBS 0.0198f
C8044 VDD.n989 VSUBS 0.0455f
C8045 VDD.n990 VSUBS 0.0842f
C8046 VDD.n991 VSUBS 0.0198f
C8047 VDD.n992 VSUBS 0.0455f
C8048 VDD.n993 VSUBS 0.0842f
C8049 VDD.n994 VSUBS 0.0198f
C8050 VDD.n995 VSUBS 0.0455f
C8051 VDD.n996 VSUBS 0.0842f
C8052 VDD.n997 VSUBS 0.0198f
C8053 VDD.n998 VSUBS 0.0455f
C8054 VDD.n999 VSUBS 0.0842f
C8055 VDD.n1000 VSUBS 0.0198f
C8056 VDD.n1001 VSUBS 0.0455f
C8057 VDD.n1002 VSUBS 0.0842f
C8058 VDD.n1003 VSUBS 0.0198f
C8059 VDD.n1004 VSUBS 0.0455f
C8060 VDD.n1005 VSUBS 0.0842f
C8061 VDD.n1006 VSUBS 0.0198f
C8062 VDD.n1007 VSUBS 0.0455f
C8063 VDD.n1008 VSUBS 0.0842f
C8064 VDD.n1009 VSUBS 0.0198f
C8065 VDD.n1010 VSUBS 0.0455f
C8066 VDD.n1011 VSUBS 0.0842f
C8067 VDD.n1012 VSUBS 0.0198f
C8068 VDD.n1013 VSUBS 0.0455f
C8069 VDD.n1014 VSUBS 0.0842f
C8070 VDD.n1015 VSUBS 0.0198f
C8071 VDD.n1016 VSUBS 0.0264f
C8072 VDD.n1017 VSUBS 0.0227f
C8073 VDD.n1018 VSUBS 0.539f
C8074 VDD.n1019 VSUBS 0.0198f
C8075 VDD.n1020 VSUBS 0.0405f
C8076 VDD.n1021 VSUBS 0.0405f
C8077 VDD.n1022 VSUBS 0.0198f
C8078 VDD.n1023 VSUBS 0.0405f
C8079 VDD.n1024 VSUBS 0.0405f
C8080 VDD.n1025 VSUBS 0.0198f
C8081 VDD.n1026 VSUBS 0.0405f
C8082 VDD.n1027 VSUBS 0.0405f
C8083 VDD.n1028 VSUBS 0.0198f
C8084 VDD.n1029 VSUBS 0.0405f
C8085 VDD.n1030 VSUBS 0.0405f
C8086 VDD.n1031 VSUBS 0.0198f
C8087 VDD.n1032 VSUBS 0.0405f
C8088 VDD.n1033 VSUBS 0.0405f
C8089 VDD.n1034 VSUBS 0.0198f
C8090 VDD.n1035 VSUBS 0.0405f
C8091 VDD.n1036 VSUBS 0.0405f
C8092 VDD.n1037 VSUBS 0.0198f
C8093 VDD.n1038 VSUBS 0.0405f
C8094 VDD.n1039 VSUBS 0.0405f
C8095 VDD.n1040 VSUBS 0.0198f
C8096 VDD.n1041 VSUBS 0.0405f
C8097 VDD.n1042 VSUBS 0.0405f
C8098 VDD.n1043 VSUBS 0.0198f
C8099 VDD.n1044 VSUBS 0.0405f
C8100 VDD.n1045 VSUBS 0.0405f
C8101 VDD.n1046 VSUBS 0.0198f
C8102 VDD.n1047 VSUBS 0.0405f
C8103 VDD.n1048 VSUBS 0.0405f
C8104 VDD.n1049 VSUBS 0.0198f
C8105 VDD.n1050 VSUBS 0.0405f
C8106 VDD.n1051 VSUBS 0.0405f
C8107 VDD.n1052 VSUBS 0.0198f
C8108 VDD.n1053 VSUBS 0.0405f
C8109 VDD.n1054 VSUBS 0.0405f
C8110 VDD.n1055 VSUBS 0.0198f
C8111 VDD.n1056 VSUBS 0.0405f
C8112 VDD.n1057 VSUBS 0.0155f
C8113 VDD.n1058 VSUBS 0.0405f
C8114 VDD.n1059 VSUBS 0.0198f
C8115 VDD.n1060 VSUBS 0.0405f
C8116 VDD.n1061 VSUBS 0.0155f
C8117 VDD.n1062 VSUBS 0.0405f
C8118 VDD.n1063 VSUBS 0.0198f
C8119 VDD.n1064 VSUBS 0.0405f
C8120 VDD.n1065 VSUBS 0.0155f
C8121 VDD.n1066 VSUBS 0.0405f
C8122 VDD.n1067 VSUBS 0.0198f
C8123 VDD.n1068 VSUBS 0.0405f
C8124 VDD.n1069 VSUBS 0.0155f
C8125 VDD.n1070 VSUBS 0.0405f
C8126 VDD.n1071 VSUBS 0.0198f
C8127 VDD.n1072 VSUBS 0.0405f
C8128 VDD.n1073 VSUBS 0.0155f
C8129 VDD.n1074 VSUBS 0.0405f
C8130 VDD.n1075 VSUBS 0.0198f
C8131 VDD.n1076 VSUBS 0.0405f
C8132 VDD.n1077 VSUBS 0.0327f
C8133 VDD.n1078 VSUBS 0.0405f
C8134 VDD.n1079 VSUBS 0.0198f
C8135 VDD.n1080 VSUBS 0.0614f
C8136 VDD.n1081 VSUBS 0.0842f
C8137 VDD.n1082 VSUBS 0.0198f
C8138 VDD.n1083 VSUBS 0.0842f
C8139 VDD.n1084 VSUBS 0.0198f
C8140 VDD.n1086 VSUBS 0.0595f
C8141 VDD.n1087 VSUBS 0.0198f
C8142 VDD.n1088 VSUBS 0.00989f
C8143 VDD.n1089 VSUBS 0.00989f
C8144 VDD.n1090 VSUBS 0.0842f
C8145 VDD.n1091 VSUBS 0.0198f
C8146 VDD.n1092 VSUBS 0.0842f
C8147 VDD.n1093 VSUBS 0.0198f
C8148 VDD.n1095 VSUBS 0.0198f
C8149 VDD.n1096 VSUBS 0.0842f
C8150 VDD.n1097 VSUBS 0.0198f
C8151 VDD.n1098 VSUBS 0.0842f
C8152 VDD.n1099 VSUBS 0.0198f
C8153 VDD.n1101 VSUBS 0.0842f
C8154 VDD.n1102 VSUBS 0.0198f
C8155 VDD.n1103 VSUBS 0.207f
C8156 VDD.n1104 VSUBS 0.237f
C8157 VDD.n1105 VSUBS 0.0842f
C8158 VDD.n1106 VSUBS 0.0198f
C8159 VDD.n1107 VSUBS 0.0455f
C8160 VDD.n1108 VSUBS 0.0842f
C8161 VDD.n1109 VSUBS 0.0198f
C8162 VDD.n1110 VSUBS 0.0455f
C8163 VDD.n1111 VSUBS 0.0842f
C8164 VDD.n1112 VSUBS 0.0198f
C8165 VDD.n1113 VSUBS 0.0455f
C8166 VDD.n1114 VSUBS 0.0842f
C8167 VDD.n1115 VSUBS 0.0198f
C8168 VDD.n1116 VSUBS 0.0455f
C8169 VDD.n1117 VSUBS 0.0842f
C8170 VDD.n1118 VSUBS 0.0198f
C8171 VDD.n1119 VSUBS 0.0455f
C8172 VDD.n1120 VSUBS 0.0842f
C8173 VDD.n1121 VSUBS 0.0198f
C8174 VDD.n1122 VSUBS 0.0455f
C8175 VDD.n1123 VSUBS 0.0842f
C8176 VDD.n1124 VSUBS 0.0198f
C8177 VDD.n1125 VSUBS 0.0455f
C8178 VDD.n1126 VSUBS 0.0842f
C8179 VDD.n1127 VSUBS 0.0198f
C8180 VDD.n1128 VSUBS 0.0455f
C8181 VDD.n1129 VSUBS 0.0842f
C8182 VDD.n1130 VSUBS 0.0198f
C8183 VDD.n1131 VSUBS 0.0455f
C8184 VDD.n1132 VSUBS 0.0842f
C8185 VDD.n1133 VSUBS 0.0198f
C8186 VDD.n1134 VSUBS 0.0455f
C8187 VDD.n1135 VSUBS 0.0842f
C8188 VDD.n1136 VSUBS 0.0198f
C8189 VDD.n1137 VSUBS 0.0455f
C8190 VDD.n1138 VSUBS 0.0842f
C8191 VDD.n1139 VSUBS 0.0198f
C8192 VDD.n1140 VSUBS 0.0455f
C8193 VDD.n1141 VSUBS 0.0842f
C8194 VDD.n1142 VSUBS 0.0198f
C8195 VDD.n1143 VSUBS 0.0455f
C8196 VDD.n1144 VSUBS 0.0842f
C8197 VDD.n1145 VSUBS 0.0198f
C8198 VDD.n1146 VSUBS 0.0455f
C8199 VDD.n1147 VSUBS 0.0842f
C8200 VDD.n1148 VSUBS 0.0198f
C8201 VDD.n1149 VSUBS 0.0455f
C8202 VDD.n1150 VSUBS 0.0842f
C8203 VDD.n1151 VSUBS 0.0198f
C8204 VDD.n1152 VSUBS 0.0455f
C8205 VDD.n1153 VSUBS 0.0842f
C8206 VDD.n1154 VSUBS 0.0198f
C8207 VDD.n1155 VSUBS 0.0441f
C8208 VDD.n1156 VSUBS 0.0842f
C8209 VDD.n1157 VSUBS 0.0198f
C8210 VDD.n1158 VSUBS 0.0909f
C8211 VDD.n1159 VSUBS 0.0842f
C8212 VDD.n1160 VSUBS 0.0198f
C8213 VDD.n1161 VSUBS 0.0955f
C8214 VDD.n1162 VSUBS 0.0842f
C8215 VDD.n1163 VSUBS 0.0198f
C8216 VDD.n1164 VSUBS 0.0955f
C8217 VDD.n1165 VSUBS 0.0842f
C8218 VDD.n1166 VSUBS 0.0198f
C8219 VDD.n1167 VSUBS 0.0955f
C8220 VDD.n1168 VSUBS 0.0842f
C8221 VDD.n1169 VSUBS 0.0198f
C8222 VDD.n1170 VSUBS 0.0955f
C8223 VDD.n1171 VSUBS 0.0842f
C8224 VDD.n1172 VSUBS 0.0198f
C8225 VDD.n1173 VSUBS 0.0955f
C8226 VDD.n1174 VSUBS 0.0842f
C8227 VDD.n1175 VSUBS 0.0198f
C8228 VDD.n1176 VSUBS 0.0955f
C8229 VDD.n1177 VSUBS 0.0842f
C8230 VDD.n1178 VSUBS 0.0198f
C8231 VDD.n1179 VSUBS 0.0955f
C8232 VDD.n1180 VSUBS 0.0842f
C8233 VDD.n1181 VSUBS 0.0198f
C8234 VDD.n1182 VSUBS 0.0955f
C8235 VDD.n1183 VSUBS 0.0842f
C8236 VDD.n1184 VSUBS 0.0198f
C8237 VDD.n1185 VSUBS 0.0955f
C8238 VDD.n1186 VSUBS 0.0842f
C8239 VDD.n1187 VSUBS 0.0198f
C8240 VDD.n1188 VSUBS 0.0899f
C8241 VDD.n1189 VSUBS 0.327f
C8242 VDD.n1190 VSUBS 0.0325f
C8243 VDD.n1191 VSUBS 0.335f
C8244 VDD.n1192 VSUBS 0.0155f
C8245 VDD.n1193 VSUBS 0.135f
C8246 VDD.n1194 VSUBS 0.0155f
C8247 VDD.n1195 VSUBS 0.167f
C8248 VDD.n1196 VSUBS 0.0155f
C8249 VDD.n1197 VSUBS 0.167f
C8250 VDD.n1198 VSUBS 0.0155f
C8251 VDD.n1199 VSUBS 0.167f
C8252 VDD.n1200 VSUBS 0.0155f
C8253 VDD.n1201 VSUBS 0.167f
C8254 VDD.n1202 VSUBS 0.0155f
C8255 VDD.n1203 VSUBS 0.167f
C8256 VDD.n1204 VSUBS 0.0155f
C8257 VDD.n1205 VSUBS 0.115f
C8258 VDD.n1206 VSUBS 0.385f
C8259 VDD.n1207 VSUBS 2.82f
C8260 VDD.n1208 VSUBS 1.76f
C8261 VDD.t38 VSUBS 0.0114f
C8262 VDD.t40 VSUBS 0.0114f
C8263 VDD.n1209 VSUBS 0.0411f
C8264 VDD.n1210 VSUBS 0.0155f
C8265 VDD.n1211 VSUBS 0.167f
C8266 VDD.n1212 VSUBS 0.0155f
C8267 VDD.n1213 VSUBS 0.167f
C8268 VDD.n1214 VSUBS 0.0155f
C8269 VDD.n1215 VSUBS 0.167f
C8270 VDD.n1216 VSUBS 0.0155f
C8271 VDD.n1217 VSUBS 0.167f
C8272 VDD.n1218 VSUBS 0.0155f
C8273 VDD.n1219 VSUBS 0.167f
C8274 VDD.n1220 VSUBS 0.0155f
C8275 VDD.n1221 VSUBS 0.092f
C8276 VDD.n1222 VSUBS 0.0155f
C8277 VDD.n1223 VSUBS 0.00909f
C8278 VDD.n1225 VSUBS 0.0155f
C8279 VDD.n1226 VSUBS 0.00909f
C8280 VDD.n1227 VSUBS 0.0155f
C8281 VDD.n1228 VSUBS 0.00909f
C8282 VDD.n1229 VSUBS 0.0343f
C8283 VDD.n1231 VSUBS 0.332f
C8284 VDD.n1233 VSUBS 0.0155f
C8285 VDD.n1234 VSUBS 0.00989f
C8286 VDD.n1235 VSUBS 0.0356f
C8287 VDD.n1236 VSUBS 0.0155f
C8288 VDD.n1237 VSUBS 0.00989f
C8289 VDD.n1238 VSUBS 0.0155f
C8290 VDD.n1239 VSUBS 0.00909f
C8291 VDD.n1240 VSUBS 0.0155f
C8292 VDD.n1241 VSUBS 0.00909f
C8293 VDD.n1243 VSUBS 0.0155f
C8294 VDD.n1244 VSUBS 0.00909f
C8295 VDD.n1245 VSUBS 0.0155f
C8296 VDD.n1246 VSUBS 0.00909f
C8297 VDD.n1247 VSUBS 0.0356f
C8298 VDD.n1249 VSUBS 0.347f
C8299 VDD.n1251 VSUBS 0.0155f
C8300 VDD.n1252 VSUBS 0.00989f
C8301 VDD.n1253 VSUBS 0.0155f
C8302 VDD.n1254 VSUBS 0.0859f
C8303 VDD.n1255 VSUBS 0.0888f
C8304 VDD.n1256 VSUBS 0.0155f
C8305 VDD.n1257 VSUBS 0.15f
C8306 VDD.n1258 VSUBS 0.27f
C8307 VDD.n1259 VSUBS 0.0217f
C8308 VDD.n1260 VSUBS 0.0834f
C8309 VDD.n1261 VSUBS 0.0155f
C8310 VDD.n1262 VSUBS 0.0834f
C8311 VDD.t39 VSUBS 0.0968f
C8312 VDD.n1263 VSUBS 0.13f
C8313 VDD.n1264 VSUBS 0.0155f
C8314 VDD.n1265 VSUBS 0.0834f
C8315 VDD.n1266 VSUBS 0.0155f
C8316 VDD.n1267 VSUBS 0.0834f
C8317 VDD.n1268 VSUBS 0.161f
C8318 VDD.n1269 VSUBS 0.0155f
C8319 VDD.n1270 VSUBS 0.0834f
C8320 VDD.n1271 VSUBS 0.0155f
C8321 VDD.n1272 VSUBS 0.0834f
C8322 VDD.n1273 VSUBS 0.161f
C8323 VDD.n1274 VSUBS 0.0155f
C8324 VDD.n1275 VSUBS 0.0834f
C8325 VDD.n1276 VSUBS 0.0155f
C8326 VDD.n1277 VSUBS 0.0834f
C8327 VDD.t37 VSUBS 0.0968f
C8328 VDD.n1278 VSUBS 0.13f
C8329 VDD.n1279 VSUBS 0.0155f
C8330 VDD.n1280 VSUBS 0.0834f
C8331 VDD.n1281 VSUBS 0.0155f
C8332 VDD.n1282 VSUBS 0.0834f
C8333 VDD.n1283 VSUBS 0.27f
C8334 VDD.n1284 VSUBS 0.0217f
C8335 VDD.n1285 VSUBS 0.0834f
C8336 VDD.n1286 VSUBS 0.0155f
C8337 VDD.n1287 VSUBS 0.0982f
C8338 VDD.n1288 VSUBS 0.0155f
C8339 VDD.n1289 VSUBS 0.135f
C8340 VDD.n1290 VSUBS 0.0888f
C8341 VDD.n1291 VSUBS 0.0155f
C8342 VDD.n1292 VSUBS 0.115f
C8343 VDD.n1293 VSUBS 0.0155f
C8344 VDD.n1294 VSUBS 0.104f
C8345 VDD.n1295 VSUBS 0.255f
C8346 VDD.n1296 VSUBS 0.0204f
C8347 VDD.n1297 VSUBS 0.0834f
C8348 VDD.n1298 VSUBS 0.0155f
C8349 VDD.n1299 VSUBS 0.0834f
C8350 VDD.n1300 VSUBS 0.145f
C8351 VDD.n1301 VSUBS 0.0155f
C8352 VDD.n1302 VSUBS 0.0834f
C8353 VDD.n1303 VSUBS 0.0155f
C8354 VDD.n1304 VSUBS 0.0834f
C8355 VDD.t35 VSUBS 0.0968f
C8356 VDD.n1305 VSUBS 0.145f
C8357 VDD.n1306 VSUBS 0.0155f
C8358 VDD.n1307 VSUBS 0.0834f
C8359 VDD.n1308 VSUBS 0.0155f
C8360 VDD.n1309 VSUBS 0.0834f
C8361 VDD.n1310 VSUBS 0.255f
C8362 VDD.n1311 VSUBS 0.0307f
C8363 VDD.n1312 VSUBS 0.0834f
C8364 VDD.n1313 VSUBS 0.0155f
C8365 VDD.n1314 VSUBS 0.113f
C8366 VDD.n1315 VSUBS 0.0834f
C8367 VDD.n1316 VSUBS 0.0155f
C8368 VDD.n1317 VSUBS 0.117f
C8369 VDD.n1318 VSUBS 0.0155f
C8370 VDD.n1319 VSUBS 0.158f
C8371 VDD.n1320 VSUBS 0.0853f
C8372 VDD.n1321 VSUBS 0.0155f
C8373 VDD.n1322 VSUBS 0.00909f
C8374 VDD.n1323 VSUBS 0.0343f
C8375 VDD.n1324 VSUBS 0.0155f
C8376 VDD.n1325 VSUBS 0.00989f
C8377 VDD.n1326 VSUBS 0.0243f
C8378 VDD.n1327 VSUBS 0.0243f
C8379 VDD.n1328 VSUBS 0.0155f
C8380 VDD.n1329 VSUBS 0.0243f
C8381 VDD.n1330 VSUBS 0.0155f
C8382 VDD.n1331 VSUBS 0.0243f
C8383 VDD.n1332 VSUBS 0.0217f
C8384 VDD.n1333 VSUBS 0.034f
C8385 VDD.n1334 VSUBS 0.049f
C8386 VDD.n1335 VSUBS 0.0217f
C8387 VDD.n1336 VSUBS 0.034f
C8388 VDD.n1337 VSUBS 0.0155f
C8389 VDD.n1338 VSUBS 0.0243f
C8390 VDD.n1339 VSUBS 0.0155f
C8391 VDD.n1340 VSUBS 0.0243f
C8392 VDD.n1341 VSUBS 0.0155f
C8393 VDD.n1342 VSUBS 0.0243f
C8394 VDD.n1343 VSUBS 0.0155f
C8395 VDD.n1344 VSUBS 0.0243f
C8396 VDD.n1345 VSUBS 0.0217f
C8397 VDD.n1346 VSUBS 0.034f
C8398 VDD.n1347 VSUBS 0.047f
C8399 VDD.n1348 VSUBS 0.0204f
C8400 VDD.n1349 VSUBS 0.032f
C8401 VDD.n1350 VSUBS 0.0155f
C8402 VDD.n1351 VSUBS 0.0243f
C8403 VDD.n1352 VSUBS 0.0155f
C8404 VDD.n1353 VSUBS 0.0243f
C8405 VDD.n1354 VSUBS 0.0307f
C8406 VDD.n1355 VSUBS 0.0709f
C8407 VDD.n1356 VSUBS 0.0323f
C8408 VDD.n1357 VSUBS 0.223f
C8409 VDD.n1359 VSUBS 0.0155f
C8410 VDD.n1360 VSUBS 0.0824f
C8411 VDD.n1361 VSUBS 0.0155f
C8412 VDD.n1362 VSUBS 0.0824f
C8413 VDD.n1364 VSUBS 0.0155f
C8414 VDD.n1365 VSUBS 0.0824f
C8415 VDD.n1366 VSUBS 0.0155f
C8416 VDD.n1367 VSUBS 0.0824f
C8417 VDD.n1368 VSUBS 0.429f
C8418 VDD.n1370 VSUBS 0.0323f
C8419 VDD.n1371 VSUBS 0.0878f
C8420 VDD.n1372 VSUBS 0.561f
C8421 VDD.n1373 VSUBS 0.63f
C8422 VDD.n1374 VSUBS 1.47f
C8423 VDD.t160 VSUBS 0.0114f
C8424 VDD.t162 VSUBS 0.0114f
C8425 VDD.n1375 VSUBS 0.0413f
C8426 VDD.t156 VSUBS 0.0114f
C8427 VDD.t158 VSUBS 0.0114f
C8428 VDD.n1376 VSUBS 0.0414f
C8429 VDD.t60 VSUBS 0.0114f
C8430 VDD.t58 VSUBS 0.0114f
C8431 VDD.n1377 VSUBS 0.0413f
C8432 VDD.t54 VSUBS 0.0114f
C8433 VDD.t56 VSUBS 0.0114f
C8434 VDD.n1378 VSUBS 0.0413f
C8435 VDD.n1379 VSUBS 0.0356f
C8436 VDD.n1380 VSUBS 0.0155f
C8437 VDD.n1381 VSUBS 0.00989f
C8438 VDD.n1382 VSUBS 0.0243f
C8439 VDD.n1383 VSUBS 0.0243f
C8440 VDD.n1384 VSUBS 0.0243f
C8441 VDD.n1385 VSUBS 0.0217f
C8442 VDD.n1386 VSUBS 0.034f
C8443 VDD.n1387 VSUBS 0.049f
C8444 VDD.n1388 VSUBS 0.0217f
C8445 VDD.n1389 VSUBS 0.034f
C8446 VDD.n1390 VSUBS 0.0155f
C8447 VDD.n1391 VSUBS 0.0243f
C8448 VDD.n1392 VSUBS 0.0155f
C8449 VDD.n1393 VSUBS 0.0243f
C8450 VDD.n1394 VSUBS 0.0155f
C8451 VDD.n1395 VSUBS 0.0243f
C8452 VDD.n1396 VSUBS 0.0155f
C8453 VDD.n1397 VSUBS 0.0243f
C8454 VDD.n1398 VSUBS 0.0217f
C8455 VDD.n1399 VSUBS 0.034f
C8456 VDD.n1400 VSUBS 0.049f
C8457 VDD.n1401 VSUBS 0.0217f
C8458 VDD.n1402 VSUBS 0.034f
C8459 VDD.n1403 VSUBS 0.0155f
C8460 VDD.n1404 VSUBS 0.0243f
C8461 VDD.n1405 VSUBS 0.0155f
C8462 VDD.n1406 VSUBS 0.0243f
C8463 VDD.n1407 VSUBS 0.0155f
C8464 VDD.n1408 VSUBS 0.0243f
C8465 VDD.n1409 VSUBS 0.0155f
C8466 VDD.n1410 VSUBS 0.0243f
C8467 VDD.n1411 VSUBS 0.0318f
C8468 VDD.n1412 VSUBS 0.0703f
C8469 VDD.n1413 VSUBS 0.0337f
C8470 VDD.n1414 VSUBS 0.235f
C8471 VDD.n1416 VSUBS 0.0155f
C8472 VDD.n1417 VSUBS 0.0848f
C8473 VDD.n1418 VSUBS 0.0155f
C8474 VDD.n1419 VSUBS 0.0848f
C8475 VDD.n1421 VSUBS 0.0155f
C8476 VDD.n1422 VSUBS 0.0848f
C8477 VDD.n1423 VSUBS 0.0155f
C8478 VDD.n1424 VSUBS 0.0848f
C8479 VDD.n1425 VSUBS 0.444f
C8480 VDD.n1427 VSUBS 0.0337f
C8481 VDD.n1428 VSUBS 0.0923f
C8482 VDD.n1429 VSUBS 0.0155f
C8483 VDD.n1430 VSUBS 0.00909f
C8484 VDD.n1432 VSUBS 0.0155f
C8485 VDD.n1433 VSUBS 0.00909f
C8486 VDD.n1435 VSUBS 0.0155f
C8487 VDD.n1436 VSUBS 0.00909f
C8488 VDD.n1438 VSUBS 0.0155f
C8489 VDD.n1439 VSUBS 0.00909f
C8490 VDD.n1440 VSUBS 0.0356f
C8491 VDD.n1442 VSUBS 0.347f
C8492 VDD.n1444 VSUBS 0.0155f
C8493 VDD.n1445 VSUBS 0.00989f
C8494 VDD.n1446 VSUBS 0.0155f
C8495 VDD.n1447 VSUBS 0.0834f
C8496 VDD.t59 VSUBS 0.0968f
C8497 VDD.n1448 VSUBS 0.13f
C8498 VDD.n1449 VSUBS 0.0155f
C8499 VDD.n1450 VSUBS 0.0834f
C8500 VDD.n1451 VSUBS 0.0155f
C8501 VDD.n1452 VSUBS 0.0834f
C8502 VDD.n1453 VSUBS 0.161f
C8503 VDD.n1454 VSUBS 0.0155f
C8504 VDD.n1455 VSUBS 0.0834f
C8505 VDD.n1456 VSUBS 0.0155f
C8506 VDD.n1457 VSUBS 0.0834f
C8507 VDD.n1458 VSUBS 0.161f
C8508 VDD.n1459 VSUBS 0.0155f
C8509 VDD.n1460 VSUBS 0.0834f
C8510 VDD.n1461 VSUBS 0.0155f
C8511 VDD.n1462 VSUBS 0.0834f
C8512 VDD.t57 VSUBS 0.0968f
C8513 VDD.n1463 VSUBS 0.13f
C8514 VDD.n1464 VSUBS 0.0155f
C8515 VDD.n1465 VSUBS 0.0834f
C8516 VDD.n1466 VSUBS 0.0155f
C8517 VDD.n1467 VSUBS 0.0834f
C8518 VDD.n1468 VSUBS 0.27f
C8519 VDD.n1469 VSUBS 0.0217f
C8520 VDD.n1470 VSUBS 0.0834f
C8521 VDD.n1471 VSUBS 0.0155f
C8522 VDD.n1472 VSUBS 0.15f
C8523 VDD.n1473 VSUBS 0.0888f
C8524 VDD.n1474 VSUBS 0.0155f
C8525 VDD.n1475 VSUBS 0.0908f
C8526 VDD.n1476 VSUBS 0.0155f
C8527 VDD.n1477 VSUBS 0.142f
C8528 VDD.n1478 VSUBS 0.27f
C8529 VDD.n1479 VSUBS 0.0217f
C8530 VDD.n1480 VSUBS 0.0834f
C8531 VDD.n1481 VSUBS 0.0155f
C8532 VDD.n1482 VSUBS 0.0834f
C8533 VDD.t53 VSUBS 0.0968f
C8534 VDD.n1483 VSUBS 0.13f
C8535 VDD.n1484 VSUBS 0.0155f
C8536 VDD.n1485 VSUBS 0.0834f
C8537 VDD.n1486 VSUBS 0.0155f
C8538 VDD.n1487 VSUBS 0.0834f
C8539 VDD.n1488 VSUBS 0.161f
C8540 VDD.n1489 VSUBS 0.0155f
C8541 VDD.n1490 VSUBS 0.0834f
C8542 VDD.n1491 VSUBS 0.0155f
C8543 VDD.n1492 VSUBS 0.0834f
C8544 VDD.n1493 VSUBS 0.161f
C8545 VDD.n1494 VSUBS 0.0155f
C8546 VDD.n1495 VSUBS 0.0834f
C8547 VDD.n1496 VSUBS 0.0155f
C8548 VDD.n1497 VSUBS 0.0834f
C8549 VDD.t55 VSUBS 0.0968f
C8550 VDD.n1498 VSUBS 0.13f
C8551 VDD.n1499 VSUBS 0.0155f
C8552 VDD.n1500 VSUBS 0.0834f
C8553 VDD.n1501 VSUBS 0.0155f
C8554 VDD.n1502 VSUBS 0.0834f
C8555 VDD.n1503 VSUBS 0.27f
C8556 VDD.n1504 VSUBS 0.0318f
C8557 VDD.n1505 VSUBS 0.0834f
C8558 VDD.n1506 VSUBS 0.0155f
C8559 VDD.n1507 VSUBS 0.108f
C8560 VDD.n1508 VSUBS 0.0155f
C8561 VDD.n1509 VSUBS 0.11f
C8562 VDD.n1510 VSUBS 0.0834f
C8563 VDD.n1511 VSUBS 0.0155f
C8564 VDD.n1512 VSUBS 0.14f
C8565 VDD.n1513 VSUBS 0.0155f
C8566 VDD.n1514 VSUBS 0.133f
C8567 VDD.n1515 VSUBS 0.108f
C8568 VDD.n1516 VSUBS 0.0155f
C8569 VDD.n1517 VSUBS 0.0155f
C8570 VDD.n1518 VSUBS 0.164f
C8571 VDD.n1519 VSUBS 0.165f
C8572 VDD.n1520 VSUBS 0.0155f
C8573 VDD.n1521 VSUBS 0.167f
C8574 VDD.n1522 VSUBS 0.0155f
C8575 VDD.n1523 VSUBS 0.109f
C8576 VDD.n1524 VSUBS 0.581f
C8577 VDD.n1525 VSUBS 0.408f
C8578 VDD.n1526 VSUBS 0.671f
C8579 VDD.n1527 VSUBS 0.831f
C8580 VDD.n1528 VSUBS 0.83f
C8581 VDD.n1529 VSUBS 0.628f
C8582 VDD.n1530 VSUBS 0.0243f
C8583 VDD.n1531 VSUBS 0.0243f
C8584 VDD.n1532 VSUBS 0.034f
C8585 VDD.n1533 VSUBS 0.0243f
C8586 VDD.n1534 VSUBS 0.034f
C8587 VDD.n1535 VSUBS 0.049f
C8588 VDD.n1536 VSUBS 0.0356f
C8589 VDD.n1537 VSUBS 0.0155f
C8590 VDD.n1538 VSUBS 0.00989f
C8591 VDD.n1539 VSUBS 0.0155f
C8592 VDD.n1540 VSUBS 0.00909f
C8593 VDD.n1541 VSUBS 0.0155f
C8594 VDD.n1542 VSUBS 0.00909f
C8595 VDD.n1544 VSUBS 0.0155f
C8596 VDD.n1545 VSUBS 0.00909f
C8597 VDD.n1546 VSUBS 0.0155f
C8598 VDD.n1547 VSUBS 0.00909f
C8599 VDD.n1548 VSUBS 0.0356f
C8600 VDD.n1550 VSUBS 0.347f
C8601 VDD.n1552 VSUBS 0.0155f
C8602 VDD.n1553 VSUBS 0.00989f
C8603 VDD.n1554 VSUBS 0.0356f
C8604 VDD.n1555 VSUBS 0.0155f
C8605 VDD.n1556 VSUBS 0.00989f
C8606 VDD.n1557 VSUBS 0.0155f
C8607 VDD.n1558 VSUBS 0.00909f
C8608 VDD.n1559 VSUBS 0.0155f
C8609 VDD.n1560 VSUBS 0.00909f
C8610 VDD.n1562 VSUBS 0.0155f
C8611 VDD.n1563 VSUBS 0.00909f
C8612 VDD.n1564 VSUBS 0.0155f
C8613 VDD.n1565 VSUBS 0.00909f
C8614 VDD.n1566 VSUBS 0.0356f
C8615 VDD.n1568 VSUBS 0.347f
C8616 VDD.n1570 VSUBS 0.0155f
C8617 VDD.n1571 VSUBS 0.00989f
C8618 VDD.n1572 VSUBS 0.27f
C8619 VDD.n1573 VSUBS 0.0217f
C8620 VDD.n1574 VSUBS 0.0834f
C8621 VDD.n1575 VSUBS 0.0155f
C8622 VDD.n1576 VSUBS 0.0933f
C8623 VDD.n1577 VSUBS 0.0155f
C8624 VDD.n1578 VSUBS 0.14f
C8625 VDD.n1579 VSUBS 0.0888f
C8626 VDD.n1580 VSUBS 0.0155f
C8627 VDD.n1581 VSUBS 0.11f
C8628 VDD.n1582 VSUBS 0.0155f
C8629 VDD.n1583 VSUBS 0.123f
C8630 VDD.n1584 VSUBS 0.27f
C8631 VDD.n1585 VSUBS 0.0217f
C8632 VDD.n1586 VSUBS 0.0834f
C8633 VDD.n1587 VSUBS 0.0155f
C8634 VDD.n1588 VSUBS 0.0834f
C8635 VDD.t157 VSUBS 0.0968f
C8636 VDD.n1589 VSUBS 0.0155f
C8637 VDD.n1590 VSUBS 0.13f
C8638 VDD.n1591 VSUBS 0.0155f
C8639 VDD.n1592 VSUBS 0.0834f
C8640 VDD.n1593 VSUBS 0.0155f
C8641 VDD.n1594 VSUBS 0.0834f
C8642 VDD.n1595 VSUBS 0.0155f
C8643 VDD.n1596 VSUBS 0.161f
C8644 VDD.n1597 VSUBS 0.0155f
C8645 VDD.n1598 VSUBS 0.0834f
C8646 VDD.n1599 VSUBS 0.0155f
C8647 VDD.n1600 VSUBS 0.0834f
C8648 VDD.n1601 VSUBS 0.0155f
C8649 VDD.n1602 VSUBS 0.161f
C8650 VDD.n1603 VSUBS 0.0155f
C8651 VDD.n1604 VSUBS 0.0834f
C8652 VDD.n1605 VSUBS 0.0155f
C8653 VDD.n1606 VSUBS 0.0834f
C8654 VDD.t155 VSUBS 0.0968f
C8655 VDD.n1607 VSUBS 0.0155f
C8656 VDD.n1608 VSUBS 0.13f
C8657 VDD.n1609 VSUBS 0.0155f
C8658 VDD.n1610 VSUBS 0.0834f
C8659 VDD.n1611 VSUBS 0.0155f
C8660 VDD.n1612 VSUBS 0.0834f
C8661 VDD.n1613 VSUBS 0.0217f
C8662 VDD.n1614 VSUBS 0.27f
C8663 VDD.n1615 VSUBS 0.0217f
C8664 VDD.n1616 VSUBS 0.0834f
C8665 VDD.n1617 VSUBS 0.0155f
C8666 VDD.n1618 VSUBS 0.128f
C8667 VDD.n1619 VSUBS 0.0155f
C8668 VDD.n1620 VSUBS 0.106f
C8669 VDD.n1621 VSUBS 0.0888f
C8670 VDD.n1622 VSUBS 0.0155f
C8671 VDD.n1623 VSUBS 0.145f
C8672 VDD.n1624 VSUBS 0.0155f
C8673 VDD.n1625 VSUBS 0.0883f
C8674 VDD.n1626 VSUBS 0.0217f
C8675 VDD.n1627 VSUBS 0.27f
C8676 VDD.n1628 VSUBS 0.0217f
C8677 VDD.n1629 VSUBS 0.0834f
C8678 VDD.n1630 VSUBS 0.0155f
C8679 VDD.n1631 VSUBS 0.0834f
C8680 VDD.t161 VSUBS 0.0968f
C8681 VDD.n1632 VSUBS 0.0155f
C8682 VDD.n1633 VSUBS 0.13f
C8683 VDD.n1634 VSUBS 0.0155f
C8684 VDD.n1635 VSUBS 0.0834f
C8685 VDD.n1636 VSUBS 0.0155f
C8686 VDD.n1637 VSUBS 0.0834f
C8687 VDD.n1638 VSUBS 0.0155f
C8688 VDD.n1639 VSUBS 0.161f
C8689 VDD.n1640 VSUBS 0.0155f
C8690 VDD.n1641 VSUBS 0.0834f
C8691 VDD.n1642 VSUBS 0.0155f
C8692 VDD.n1643 VSUBS 0.0834f
C8693 VDD.n1644 VSUBS 0.0155f
C8694 VDD.n1645 VSUBS 0.161f
C8695 VDD.n1646 VSUBS 0.0155f
C8696 VDD.n1647 VSUBS 0.0834f
C8697 VDD.n1648 VSUBS 0.0155f
C8698 VDD.n1649 VSUBS 0.0834f
C8699 VDD.t159 VSUBS 0.0968f
C8700 VDD.n1650 VSUBS 0.0155f
C8701 VDD.n1651 VSUBS 0.13f
C8702 VDD.n1652 VSUBS 0.0155f
C8703 VDD.n1653 VSUBS 0.0834f
C8704 VDD.n1654 VSUBS 0.0155f
C8705 VDD.n1655 VSUBS 0.0834f
C8706 VDD.n1656 VSUBS 0.0217f
C8707 VDD.n1657 VSUBS 0.27f
C8708 VDD.n1658 VSUBS 0.0217f
C8709 VDD.n1659 VSUBS 0.0503f
C8710 VDD.n1660 VSUBS 0.0515f
C8711 VDD.n1661 VSUBS 0.109f
C8712 VDD.n1662 VSUBS 0.0243f
C8713 VDD.n1663 VSUBS 0.0243f
C8714 VDD.n1664 VSUBS 0.0243f
C8715 VDD.n1665 VSUBS 0.034f
C8716 VDD.n1666 VSUBS 0.0243f
C8717 VDD.n1667 VSUBS 0.0243f
C8718 VDD.n1668 VSUBS 0.034f
C8719 VDD.n1669 VSUBS 0.049f
C8720 VDD.n1670 VSUBS 0.0356f
C8721 VDD.n1671 VSUBS 0.0155f
C8722 VDD.n1672 VSUBS 0.00989f
C8723 VDD.n1673 VSUBS 0.0155f
C8724 VDD.n1674 VSUBS 0.00909f
C8725 VDD.n1675 VSUBS 0.0155f
C8726 VDD.n1676 VSUBS 0.00909f
C8727 VDD.n1678 VSUBS 0.0155f
C8728 VDD.n1679 VSUBS 0.00909f
C8729 VDD.n1680 VSUBS 0.0155f
C8730 VDD.n1681 VSUBS 0.00909f
C8731 VDD.n1682 VSUBS 0.0356f
C8732 VDD.n1684 VSUBS 0.347f
C8733 VDD.n1686 VSUBS 0.0155f
C8734 VDD.n1687 VSUBS 0.00989f
C8735 VDD.n1688 VSUBS 0.034f
C8736 VDD.n1689 VSUBS 0.0243f
C8737 VDD.n1690 VSUBS 0.034f
C8738 VDD.n1691 VSUBS 0.049f
C8739 VDD.n1692 VSUBS 0.0356f
C8740 VDD.n1693 VSUBS 0.0155f
C8741 VDD.n1694 VSUBS 0.00989f
C8742 VDD.n1695 VSUBS 0.0155f
C8743 VDD.n1696 VSUBS 0.00909f
C8744 VDD.n1697 VSUBS 0.0155f
C8745 VDD.n1698 VSUBS 0.00909f
C8746 VDD.n1700 VSUBS 0.0155f
C8747 VDD.n1701 VSUBS 0.00909f
C8748 VDD.n1702 VSUBS 0.0155f
C8749 VDD.n1703 VSUBS 0.00909f
C8750 VDD.n1704 VSUBS 0.0356f
C8751 VDD.n1706 VSUBS 0.347f
C8752 VDD.n1708 VSUBS 0.0155f
C8753 VDD.n1709 VSUBS 0.00989f
C8754 VDD.n1710 VSUBS 0.0155f
C8755 VDD.n1711 VSUBS 0.147f
C8756 VDD.n1712 VSUBS 0.27f
C8757 VDD.n1713 VSUBS 0.0217f
C8758 VDD.n1714 VSUBS 0.0834f
C8759 VDD.n1715 VSUBS 0.0155f
C8760 VDD.n1716 VSUBS 0.0834f
C8761 VDD.t446 VSUBS 0.0968f
C8762 VDD.n1717 VSUBS 0.13f
C8763 VDD.n1718 VSUBS 0.0155f
C8764 VDD.n1719 VSUBS 0.0834f
C8765 VDD.n1720 VSUBS 0.0155f
C8766 VDD.n1721 VSUBS 0.0834f
C8767 VDD.n1722 VSUBS 0.161f
C8768 VDD.n1723 VSUBS 0.0155f
C8769 VDD.n1724 VSUBS 0.0834f
C8770 VDD.n1725 VSUBS 0.0155f
C8771 VDD.n1726 VSUBS 0.0834f
C8772 VDD.n1727 VSUBS 0.0155f
C8773 VDD.n1728 VSUBS 0.161f
C8774 VDD.n1729 VSUBS 0.0155f
C8775 VDD.n1730 VSUBS 0.0834f
C8776 VDD.n1731 VSUBS 0.0155f
C8777 VDD.n1732 VSUBS 0.0834f
C8778 VDD.t452 VSUBS 0.0968f
C8779 VDD.n1733 VSUBS 0.0155f
C8780 VDD.n1734 VSUBS 0.13f
C8781 VDD.n1735 VSUBS 0.0155f
C8782 VDD.n1736 VSUBS 0.0834f
C8783 VDD.n1737 VSUBS 0.0155f
C8784 VDD.n1738 VSUBS 0.0834f
C8785 VDD.n1739 VSUBS 0.0217f
C8786 VDD.n1740 VSUBS 0.27f
C8787 VDD.n1741 VSUBS 0.0217f
C8788 VDD.n1742 VSUBS 0.0834f
C8789 VDD.n1743 VSUBS 0.0155f
C8790 VDD.n1744 VSUBS 0.103f
C8791 VDD.n1745 VSUBS 0.0155f
C8792 VDD.n1746 VSUBS 0.13f
C8793 VDD.n1747 VSUBS 0.0888f
C8794 VDD.n1748 VSUBS 0.0155f
C8795 VDD.n1749 VSUBS 0.12f
C8796 VDD.n1750 VSUBS 0.0155f
C8797 VDD.n1751 VSUBS 0.113f
C8798 VDD.n1752 VSUBS 0.0217f
C8799 VDD.n1753 VSUBS 0.27f
C8800 VDD.n1754 VSUBS 0.0217f
C8801 VDD.n1755 VSUBS 0.0834f
C8802 VDD.n1756 VSUBS 0.0155f
C8803 VDD.n1757 VSUBS 0.0834f
C8804 VDD.t31 VSUBS 0.0968f
C8805 VDD.n1758 VSUBS 0.0155f
C8806 VDD.n1759 VSUBS 0.13f
C8807 VDD.n1760 VSUBS 0.0155f
C8808 VDD.n1761 VSUBS 0.0834f
C8809 VDD.n1762 VSUBS 0.0155f
C8810 VDD.n1763 VSUBS 0.0834f
C8811 VDD.n1764 VSUBS 0.0155f
C8812 VDD.n1765 VSUBS 0.161f
C8813 VDD.n1766 VSUBS 0.0155f
C8814 VDD.n1767 VSUBS 0.0834f
C8815 VDD.n1768 VSUBS 0.0155f
C8816 VDD.n1769 VSUBS 0.0834f
C8817 VDD.n1770 VSUBS 0.0155f
C8818 VDD.n1771 VSUBS 0.161f
C8819 VDD.n1772 VSUBS 0.0155f
C8820 VDD.n1773 VSUBS 0.0834f
C8821 VDD.n1774 VSUBS 0.0155f
C8822 VDD.n1775 VSUBS 0.0834f
C8823 VDD.t140 VSUBS 0.0968f
C8824 VDD.n1776 VSUBS 0.0155f
C8825 VDD.n1777 VSUBS 0.13f
C8826 VDD.n1778 VSUBS 0.0155f
C8827 VDD.n1779 VSUBS 0.0834f
C8828 VDD.n1780 VSUBS 0.0155f
C8829 VDD.n1781 VSUBS 0.0834f
C8830 VDD.n1782 VSUBS 0.0217f
C8831 VDD.n1783 VSUBS 0.27f
C8832 VDD.n1784 VSUBS 0.0217f
C8833 VDD.n1785 VSUBS 0.0834f
C8834 VDD.n1786 VSUBS 0.0155f
C8835 VDD.n1787 VSUBS 0.137f
C8836 VDD.n1788 VSUBS 0.0155f
C8837 VDD.n1789 VSUBS 0.0957f
C8838 VDD.n1790 VSUBS 0.0888f
C8839 VDD.n1791 VSUBS 0.0155f
C8840 VDD.n1792 VSUBS 0.0982f
C8841 VDD.n1793 VSUBS 0.0331f
C8842 VDD.n1794 VSUBS 0.814f
C8843 VDD.n1795 VSUBS 2.62f
C8844 VDD.n1796 VSUBS 1.69f
C8845 VDD.n1797 VSUBS 0.00723f
C8846 VDD.n1798 VSUBS 0.00354f
C8847 VDD.n1799 VSUBS 0.0145f
C8848 VDD.t336 VSUBS 0.0114f
C8849 VDD.t283 VSUBS 0.0114f
C8850 VDD.n1800 VSUBS 0.0268f
C8851 VDD.n1801 VSUBS 0.0127f
C8852 VDD.n1802 VSUBS 0.0267f
C8853 VDD.n1803 VSUBS 0.0142f
C8854 VDD.n1804 VSUBS 0.00723f
C8855 VDD.n1805 VSUBS 0.00354f
C8856 VDD.n1806 VSUBS 0.0145f
C8857 VDD.t265 VSUBS 0.0114f
C8858 VDD.t183 VSUBS 0.0114f
C8859 VDD.n1807 VSUBS 0.0268f
C8860 VDD.n1808 VSUBS 0.0127f
C8861 VDD.n1809 VSUBS 0.0267f
C8862 VDD.n1810 VSUBS 0.0142f
C8863 VDD.n1811 VSUBS 0.00723f
C8864 VDD.n1812 VSUBS 0.00354f
C8865 VDD.n1813 VSUBS 0.0145f
C8866 VDD.t364 VSUBS 0.0114f
C8867 VDD.t316 VSUBS 0.0114f
C8868 VDD.n1814 VSUBS 0.0268f
C8869 VDD.n1815 VSUBS 0.0127f
C8870 VDD.n1816 VSUBS 0.0267f
C8871 VDD.n1817 VSUBS 0.0142f
C8872 VDD.n1818 VSUBS 0.00723f
C8873 VDD.n1819 VSUBS 0.00354f
C8874 VDD.n1820 VSUBS 0.0145f
C8875 VDD.t314 VSUBS 0.0114f
C8876 VDD.t210 VSUBS 0.0114f
C8877 VDD.n1821 VSUBS 0.0268f
C8878 VDD.n1822 VSUBS 0.0127f
C8879 VDD.n1823 VSUBS 0.0267f
C8880 VDD.n1824 VSUBS 0.0142f
C8881 VDD.n1825 VSUBS 0.00723f
C8882 VDD.n1826 VSUBS 0.00354f
C8883 VDD.n1827 VSUBS 0.0145f
C8884 VDD.t246 VSUBS 0.0114f
C8885 VDD.t213 VSUBS 0.0114f
C8886 VDD.n1828 VSUBS 0.0268f
C8887 VDD.n1829 VSUBS 0.0127f
C8888 VDD.n1830 VSUBS 0.0267f
C8889 VDD.n1831 VSUBS 0.0142f
C8890 VDD.n1832 VSUBS 0.00723f
C8891 VDD.n1833 VSUBS 0.00354f
C8892 VDD.n1834 VSUBS 0.0145f
C8893 VDD.t347 VSUBS 0.0114f
C8894 VDD.t293 VSUBS 0.0114f
C8895 VDD.n1835 VSUBS 0.0268f
C8896 VDD.n1836 VSUBS 0.0127f
C8897 VDD.n1837 VSUBS 0.0267f
C8898 VDD.n1838 VSUBS 0.0142f
C8899 VDD.n1839 VSUBS 0.00723f
C8900 VDD.n1840 VSUBS 0.00354f
C8901 VDD.n1841 VSUBS 0.0145f
C8902 VDD.t352 VSUBS 0.0114f
C8903 VDD.t192 VSUBS 0.0114f
C8904 VDD.n1842 VSUBS 0.0268f
C8905 VDD.n1843 VSUBS 0.0127f
C8906 VDD.n1844 VSUBS 0.0267f
C8907 VDD.n1845 VSUBS 0.0142f
C8908 VDD.n1846 VSUBS 0.00723f
C8909 VDD.n1847 VSUBS 0.00354f
C8910 VDD.n1848 VSUBS 0.0145f
C8911 VDD.t281 VSUBS 0.0114f
C8912 VDD.t198 VSUBS 0.0114f
C8913 VDD.n1849 VSUBS 0.0268f
C8914 VDD.n1850 VSUBS 0.0127f
C8915 VDD.n1851 VSUBS 0.0267f
C8916 VDD.n1852 VSUBS 0.0142f
C8917 VDD.n1853 VSUBS 0.00723f
C8918 VDD.n1854 VSUBS 0.00354f
C8919 VDD.n1855 VSUBS 0.0145f
C8920 VDD.t322 VSUBS 0.0114f
C8921 VDD.t273 VSUBS 0.0114f
C8922 VDD.n1856 VSUBS 0.0268f
C8923 VDD.n1857 VSUBS 0.0127f
C8924 VDD.n1858 VSUBS 0.0267f
C8925 VDD.n1859 VSUBS 0.0142f
C8926 VDD.n1860 VSUBS 0.00723f
C8927 VDD.n1861 VSUBS 0.00354f
C8928 VDD.n1862 VSUBS 0.0145f
C8929 VDD.t267 VSUBS 0.0114f
C8930 VDD.t223 VSUBS 0.0114f
C8931 VDD.n1863 VSUBS 0.0268f
C8932 VDD.n1864 VSUBS 0.0127f
C8933 VDD.n1865 VSUBS 0.0267f
C8934 VDD.n1866 VSUBS 0.0142f
C8935 VDD.n1867 VSUBS 0.00723f
C8936 VDD.n1868 VSUBS 0.00354f
C8937 VDD.n1869 VSUBS 0.0145f
C8938 VDD.t368 VSUBS 0.0114f
C8939 VDD.t174 VSUBS 0.0114f
C8940 VDD.n1870 VSUBS 0.0268f
C8941 VDD.n1871 VSUBS 0.0127f
C8942 VDD.n1872 VSUBS 0.0267f
C8943 VDD.n1873 VSUBS 0.0142f
C8944 VDD.n1874 VSUBS 0.00723f
C8945 VDD.n1875 VSUBS 0.00354f
C8946 VDD.n1876 VSUBS 0.0145f
C8947 VDD.t297 VSUBS 0.0114f
C8948 VDD.t252 VSUBS 0.0114f
C8949 VDD.n1877 VSUBS 0.0268f
C8950 VDD.n1878 VSUBS 0.0127f
C8951 VDD.n1879 VSUBS 0.0267f
C8952 VDD.n1880 VSUBS 0.0142f
C8953 VDD.n1881 VSUBS 0.00723f
C8954 VDD.n1882 VSUBS 0.00354f
C8955 VDD.n1883 VSUBS 0.0145f
C8956 VDD.t270 VSUBS 0.0114f
C8957 VDD.t351 VSUBS 0.0114f
C8958 VDD.n1884 VSUBS 0.0268f
C8959 VDD.n1885 VSUBS 0.0127f
C8960 VDD.n1886 VSUBS 0.0267f
C8961 VDD.n1887 VSUBS 0.0142f
C8962 VDD.n1888 VSUBS 0.00723f
C8963 VDD.n1889 VSUBS 0.00354f
C8964 VDD.n1890 VSUBS 0.0145f
C8965 VDD.t323 VSUBS 0.0114f
C8966 VDD.t224 VSUBS 0.0114f
C8967 VDD.n1891 VSUBS 0.0268f
C8968 VDD.n1892 VSUBS 0.0127f
C8969 VDD.n1893 VSUBS 0.0267f
C8970 VDD.n1894 VSUBS 0.0142f
C8971 VDD.n1895 VSUBS 0.00723f
C8972 VDD.n1896 VSUBS 0.00354f
C8973 VDD.n1897 VSUBS 0.0145f
C8974 VDD.t234 VSUBS 0.0114f
C8975 VDD.t274 VSUBS 0.0114f
C8976 VDD.n1898 VSUBS 0.0268f
C8977 VDD.n1899 VSUBS 0.0127f
C8978 VDD.n1900 VSUBS 0.0267f
C8979 VDD.n1901 VSUBS 0.0142f
C8980 VDD.n1902 VSUBS 0.00723f
C8981 VDD.n1903 VSUBS 0.00354f
C8982 VDD.n1904 VSUBS 0.0145f
C8983 VDD.t353 VSUBS 0.0114f
C8984 VDD.t348 VSUBS 0.0114f
C8985 VDD.n1905 VSUBS 0.0268f
C8986 VDD.n1906 VSUBS 0.0127f
C8987 VDD.n1907 VSUBS 0.0267f
C8988 VDD.n1908 VSUBS 0.0142f
C8989 VDD.n1909 VSUBS 0.00723f
C8990 VDD.n1910 VSUBS 0.00354f
C8991 VDD.n1911 VSUBS 0.0145f
C8992 VDD.t220 VSUBS 0.0114f
C8993 VDD.t253 VSUBS 0.0114f
C8994 VDD.n1912 VSUBS 0.0268f
C8995 VDD.n1913 VSUBS 0.0127f
C8996 VDD.n1914 VSUBS 0.0267f
C8997 VDD.n1915 VSUBS 0.0142f
C8998 VDD.n1916 VSUBS 0.00723f
C8999 VDD.n1917 VSUBS 0.00354f
C9000 VDD.n1918 VSUBS 0.0145f
C9001 VDD.t268 VSUBS 0.0114f
C9002 VDD.t317 VSUBS 0.0114f
C9003 VDD.n1919 VSUBS 0.0268f
C9004 VDD.n1920 VSUBS 0.0127f
C9005 VDD.n1921 VSUBS 0.0267f
C9006 VDD.n1922 VSUBS 0.0142f
C9007 VDD.n1923 VSUBS 0.00723f
C9008 VDD.n1924 VSUBS 0.00354f
C9009 VDD.n1925 VSUBS 0.0145f
C9010 VDD.t194 VSUBS 0.0114f
C9011 VDD.t277 VSUBS 0.0114f
C9012 VDD.n1926 VSUBS 0.0268f
C9013 VDD.n1927 VSUBS 0.0127f
C9014 VDD.n1928 VSUBS 0.0267f
C9015 VDD.n1929 VSUBS 0.0142f
C9016 VDD.n1930 VSUBS 0.00723f
C9017 VDD.n1931 VSUBS 0.00354f
C9018 VDD.n1932 VSUBS 0.0202f
C9019 VDD.t185 VSUBS 0.0114f
C9020 VDD.t269 VSUBS 0.0114f
C9021 VDD.n1933 VSUBS 0.0268f
C9022 VDD.n1934 VSUBS 0.0127f
C9023 VDD.n1935 VSUBS 0.0267f
C9024 VDD.n1936 VSUBS 0.0142f
C9025 VDD.n1937 VSUBS 0.215f
C9026 VDD.n1938 VSUBS 0.0867f
C9027 VDD.n1939 VSUBS 0.0867f
C9028 VDD.n1940 VSUBS 0.0867f
C9029 VDD.n1941 VSUBS 0.0867f
C9030 VDD.n1942 VSUBS 0.0867f
C9031 VDD.n1943 VSUBS 0.0867f
C9032 VDD.n1944 VSUBS 0.0867f
C9033 VDD.n1945 VSUBS 0.0867f
C9034 VDD.n1946 VSUBS 0.0867f
C9035 VDD.n1947 VSUBS 0.0867f
C9036 VDD.n1948 VSUBS 0.0867f
C9037 VDD.n1949 VSUBS 0.0867f
C9038 VDD.n1950 VSUBS 0.0867f
C9039 VDD.n1951 VSUBS 0.0867f
C9040 VDD.n1952 VSUBS 0.0867f
C9041 VDD.n1953 VSUBS 0.0867f
C9042 VDD.n1954 VSUBS 0.0867f
C9043 VDD.n1955 VSUBS 0.0867f
C9044 VDD.n1956 VSUBS 0.0867f
C9045 VDD.n1957 VSUBS 0.0867f
C9046 VDD.n1958 VSUBS 0.0867f
C9047 VDD.n1959 VSUBS 0.0867f
C9048 VDD.n1960 VSUBS 0.0867f
C9049 VDD.n1961 VSUBS 0.0867f
C9050 VDD.n1962 VSUBS 0.0867f
C9051 VDD.n1963 VSUBS 0.0867f
C9052 VDD.n1964 VSUBS 0.0867f
C9053 VDD.n1965 VSUBS 0.0867f
C9054 VDD.n1966 VSUBS 0.0867f
C9055 VDD.n1967 VSUBS 0.0867f
C9056 VDD.n1968 VSUBS 0.0867f
C9057 VDD.n1969 VSUBS 0.0867f
C9058 VDD.n1970 VSUBS 0.0867f
C9059 VDD.n1971 VSUBS 0.0867f
C9060 VDD.n1972 VSUBS 0.0867f
C9061 VDD.n1973 VSUBS 0.0867f
C9062 VDD.n1974 VSUBS 0.0867f
C9063 VDD.n1975 VSUBS 0.0867f
C9064 VDD.n1976 VSUBS 0.00717f
C9065 VDD.n1977 VSUBS 0.00349f
C9066 VDD.n1978 VSUBS 0.0145f
C9067 VDD.t349 VSUBS 0.0114f
C9068 VDD.t301 VSUBS 0.0114f
C9069 VDD.n1979 VSUBS 0.0268f
C9070 VDD.n1980 VSUBS 0.0129f
C9071 VDD.n1981 VSUBS 0.027f
C9072 VDD.n1982 VSUBS 0.0142f
C9073 VDD.n1983 VSUBS 0.00717f
C9074 VDD.n1984 VSUBS 0.00349f
C9075 VDD.n1985 VSUBS 0.0145f
C9076 VDD.t278 VSUBS 0.0114f
C9077 VDD.t196 VSUBS 0.0114f
C9078 VDD.n1986 VSUBS 0.0268f
C9079 VDD.n1987 VSUBS 0.0129f
C9080 VDD.n1988 VSUBS 0.027f
C9081 VDD.n1989 VSUBS 0.0142f
C9082 VDD.n1990 VSUBS 0.00717f
C9083 VDD.n1991 VSUBS 0.00349f
C9084 VDD.n1992 VSUBS 0.0145f
C9085 VDD.t178 VSUBS 0.0114f
C9086 VDD.t333 VSUBS 0.0114f
C9087 VDD.n1993 VSUBS 0.0268f
C9088 VDD.n1994 VSUBS 0.0129f
C9089 VDD.n1995 VSUBS 0.027f
C9090 VDD.n1996 VSUBS 0.0142f
C9091 VDD.n1997 VSUBS 0.00717f
C9092 VDD.n1998 VSUBS 0.00349f
C9093 VDD.n1999 VSUBS 0.0145f
C9094 VDD.t332 VSUBS 0.0114f
C9095 VDD.t215 VSUBS 0.0114f
C9096 VDD.n2000 VSUBS 0.0268f
C9097 VDD.n2001 VSUBS 0.0129f
C9098 VDD.n2002 VSUBS 0.027f
C9099 VDD.n2003 VSUBS 0.0142f
C9100 VDD.n2004 VSUBS 0.00717f
C9101 VDD.n2005 VSUBS 0.00349f
C9102 VDD.n2006 VSUBS 0.0145f
C9103 VDD.t260 VSUBS 0.0114f
C9104 VDD.t225 VSUBS 0.0114f
C9105 VDD.n2007 VSUBS 0.0268f
C9106 VDD.n2008 VSUBS 0.0129f
C9107 VDD.n2009 VSUBS 0.027f
C9108 VDD.n2010 VSUBS 0.0142f
C9109 VDD.n2011 VSUBS 0.00717f
C9110 VDD.n2012 VSUBS 0.00349f
C9111 VDD.n2013 VSUBS 0.0145f
C9112 VDD.t359 VSUBS 0.0114f
C9113 VDD.t311 VSUBS 0.0114f
C9114 VDD.n2014 VSUBS 0.0268f
C9115 VDD.n2015 VSUBS 0.0129f
C9116 VDD.n2016 VSUBS 0.027f
C9117 VDD.n2017 VSUBS 0.0142f
C9118 VDD.n2018 VSUBS 0.00717f
C9119 VDD.n2019 VSUBS 0.00349f
C9120 VDD.n2020 VSUBS 0.0145f
C9121 VDD.t366 VSUBS 0.0114f
C9122 VDD.t206 VSUBS 0.0114f
C9123 VDD.n2021 VSUBS 0.0268f
C9124 VDD.n2022 VSUBS 0.0129f
C9125 VDD.n2023 VSUBS 0.027f
C9126 VDD.n2024 VSUBS 0.0142f
C9127 VDD.n2025 VSUBS 0.00717f
C9128 VDD.n2026 VSUBS 0.00349f
C9129 VDD.n2027 VSUBS 0.0145f
C9130 VDD.t298 VSUBS 0.0114f
C9131 VDD.t211 VSUBS 0.0114f
C9132 VDD.n2028 VSUBS 0.0268f
C9133 VDD.n2029 VSUBS 0.0129f
C9134 VDD.n2030 VSUBS 0.027f
C9135 VDD.n2031 VSUBS 0.0142f
C9136 VDD.n2032 VSUBS 0.00717f
C9137 VDD.n2033 VSUBS 0.00349f
C9138 VDD.n2034 VSUBS 0.0145f
C9139 VDD.t339 VSUBS 0.0114f
C9140 VDD.t287 VSUBS 0.0114f
C9141 VDD.n2035 VSUBS 0.0268f
C9142 VDD.n2036 VSUBS 0.0129f
C9143 VDD.n2037 VSUBS 0.027f
C9144 VDD.n2038 VSUBS 0.0142f
C9145 VDD.n2039 VSUBS 0.00717f
C9146 VDD.n2040 VSUBS 0.00349f
C9147 VDD.n2041 VSUBS 0.0145f
C9148 VDD.t282 VSUBS 0.0114f
C9149 VDD.t230 VSUBS 0.0114f
C9150 VDD.n2042 VSUBS 0.0268f
C9151 VDD.n2043 VSUBS 0.0129f
C9152 VDD.n2044 VSUBS 0.027f
C9153 VDD.n2045 VSUBS 0.0142f
C9154 VDD.n2046 VSUBS 0.00717f
C9155 VDD.n2047 VSUBS 0.00349f
C9156 VDD.n2048 VSUBS 0.0145f
C9157 VDD.t181 VSUBS 0.0114f
C9158 VDD.t189 VSUBS 0.0114f
C9159 VDD.n2049 VSUBS 0.0268f
C9160 VDD.n2050 VSUBS 0.0129f
C9161 VDD.n2051 VSUBS 0.027f
C9162 VDD.n2052 VSUBS 0.0142f
C9163 VDD.n2053 VSUBS 0.00717f
C9164 VDD.n2054 VSUBS 0.00349f
C9165 VDD.n2055 VSUBS 0.0145f
C9166 VDD.t315 VSUBS 0.0114f
C9167 VDD.t264 VSUBS 0.0114f
C9168 VDD.n2056 VSUBS 0.0268f
C9169 VDD.n2057 VSUBS 0.0129f
C9170 VDD.n2058 VSUBS 0.027f
C9171 VDD.n2059 VSUBS 0.0142f
C9172 VDD.n2060 VSUBS 0.00717f
C9173 VDD.n2061 VSUBS 0.00349f
C9174 VDD.n2062 VSUBS 0.0145f
C9175 VDD.t286 VSUBS 0.0114f
C9176 VDD.t363 VSUBS 0.0114f
C9177 VDD.n2063 VSUBS 0.0268f
C9178 VDD.n2064 VSUBS 0.0129f
C9179 VDD.n2065 VSUBS 0.027f
C9180 VDD.n2066 VSUBS 0.0142f
C9181 VDD.n2067 VSUBS 0.00717f
C9182 VDD.n2068 VSUBS 0.00349f
C9183 VDD.n2069 VSUBS 0.0145f
C9184 VDD.t341 VSUBS 0.0114f
C9185 VDD.t231 VSUBS 0.0114f
C9186 VDD.n2070 VSUBS 0.0268f
C9187 VDD.n2071 VSUBS 0.0129f
C9188 VDD.n2072 VSUBS 0.027f
C9189 VDD.n2073 VSUBS 0.0142f
C9190 VDD.n2074 VSUBS 0.00717f
C9191 VDD.n2075 VSUBS 0.00349f
C9192 VDD.n2076 VSUBS 0.0145f
C9193 VDD.t243 VSUBS 0.0114f
C9194 VDD.t289 VSUBS 0.0114f
C9195 VDD.n2077 VSUBS 0.0268f
C9196 VDD.n2078 VSUBS 0.0129f
C9197 VDD.n2079 VSUBS 0.027f
C9198 VDD.n2080 VSUBS 0.0142f
C9199 VDD.n2081 VSUBS 0.00717f
C9200 VDD.n2082 VSUBS 0.00349f
C9201 VDD.n2083 VSUBS 0.0145f
C9202 VDD.t367 VSUBS 0.0114f
C9203 VDD.t360 VSUBS 0.0114f
C9204 VDD.n2084 VSUBS 0.0268f
C9205 VDD.n2085 VSUBS 0.0129f
C9206 VDD.n2086 VSUBS 0.027f
C9207 VDD.n2087 VSUBS 0.0142f
C9208 VDD.n2088 VSUBS 0.00717f
C9209 VDD.n2089 VSUBS 0.00349f
C9210 VDD.n2090 VSUBS 0.0145f
C9211 VDD.t228 VSUBS 0.0114f
C9212 VDD.t266 VSUBS 0.0114f
C9213 VDD.n2091 VSUBS 0.0268f
C9214 VDD.n2092 VSUBS 0.0129f
C9215 VDD.n2093 VSUBS 0.027f
C9216 VDD.n2094 VSUBS 0.0142f
C9217 VDD.n2095 VSUBS 0.00717f
C9218 VDD.n2096 VSUBS 0.00349f
C9219 VDD.n2097 VSUBS 0.0145f
C9220 VDD.t284 VSUBS 0.0114f
C9221 VDD.t338 VSUBS 0.0114f
C9222 VDD.n2098 VSUBS 0.0268f
C9223 VDD.n2099 VSUBS 0.0129f
C9224 VDD.n2100 VSUBS 0.027f
C9225 VDD.n2101 VSUBS 0.0142f
C9226 VDD.n2102 VSUBS 0.00717f
C9227 VDD.n2103 VSUBS 0.00349f
C9228 VDD.n2104 VSUBS 0.0145f
C9229 VDD.t209 VSUBS 0.0114f
C9230 VDD.t292 VSUBS 0.0114f
C9231 VDD.n2105 VSUBS 0.0268f
C9232 VDD.n2106 VSUBS 0.0129f
C9233 VDD.n2107 VSUBS 0.027f
C9234 VDD.n2108 VSUBS 0.0142f
C9235 VDD.n2109 VSUBS 0.00717f
C9236 VDD.n2110 VSUBS 0.00349f
C9237 VDD.n2111 VSUBS 0.0202f
C9238 VDD.t200 VSUBS 0.0114f
C9239 VDD.t285 VSUBS 0.0114f
C9240 VDD.n2112 VSUBS 0.0268f
C9241 VDD.n2113 VSUBS 0.0129f
C9242 VDD.n2114 VSUBS 0.027f
C9243 VDD.n2115 VSUBS 0.0142f
C9244 VDD.n2116 VSUBS 0.215f
C9245 VDD.n2117 VSUBS 0.0867f
C9246 VDD.n2118 VSUBS 0.0867f
C9247 VDD.n2119 VSUBS 0.0867f
C9248 VDD.n2120 VSUBS 0.0867f
C9249 VDD.n2121 VSUBS 0.0867f
C9250 VDD.n2122 VSUBS 0.0867f
C9251 VDD.n2123 VSUBS 0.0867f
C9252 VDD.n2124 VSUBS 0.0867f
C9253 VDD.n2125 VSUBS 0.0867f
C9254 VDD.n2126 VSUBS 0.0867f
C9255 VDD.n2127 VSUBS 0.0867f
C9256 VDD.n2128 VSUBS 0.0867f
C9257 VDD.n2129 VSUBS 0.0867f
C9258 VDD.n2130 VSUBS 0.0867f
C9259 VDD.n2131 VSUBS 0.0867f
C9260 VDD.n2132 VSUBS 0.0867f
C9261 VDD.n2133 VSUBS 0.0867f
C9262 VDD.n2134 VSUBS 0.0867f
C9263 VDD.n2135 VSUBS 0.0867f
C9264 VDD.n2136 VSUBS 0.0867f
C9265 VDD.n2137 VSUBS 0.0867f
C9266 VDD.n2138 VSUBS 0.0867f
C9267 VDD.n2139 VSUBS 0.0867f
C9268 VDD.n2140 VSUBS 0.0867f
C9269 VDD.n2141 VSUBS 0.0867f
C9270 VDD.n2142 VSUBS 0.0867f
C9271 VDD.n2143 VSUBS 0.0867f
C9272 VDD.n2144 VSUBS 0.0867f
C9273 VDD.n2145 VSUBS 0.0867f
C9274 VDD.n2146 VSUBS 0.0867f
C9275 VDD.n2147 VSUBS 0.0867f
C9276 VDD.n2148 VSUBS 0.0867f
C9277 VDD.n2149 VSUBS 0.0867f
C9278 VDD.n2150 VSUBS 0.0867f
C9279 VDD.n2151 VSUBS 0.0867f
C9280 VDD.n2152 VSUBS 0.0867f
C9281 VDD.n2153 VSUBS 0.0867f
C9282 VDD.n2154 VSUBS 0.0867f
C9283 VDD.t362 VSUBS 0.0114f
C9284 VDD.t313 VSUBS 0.0114f
C9285 VDD.n2155 VSUBS 0.0268f
C9286 VDD.n2156 VSUBS 0.0129f
C9287 VDD.n2157 VSUBS 0.00717f
C9288 VDD.n2158 VSUBS 0.00349f
C9289 VDD.n2159 VSUBS 0.0145f
C9290 VDD.n2160 VSUBS 0.0273f
C9291 VDD.n2161 VSUBS 0.0142f
C9292 VDD.t291 VSUBS 0.0114f
C9293 VDD.t208 VSUBS 0.0114f
C9294 VDD.n2162 VSUBS 0.0268f
C9295 VDD.n2163 VSUBS 0.0129f
C9296 VDD.n2164 VSUBS 0.00717f
C9297 VDD.n2165 VSUBS 0.00349f
C9298 VDD.n2166 VSUBS 0.0145f
C9299 VDD.n2167 VSUBS 0.0273f
C9300 VDD.n2168 VSUBS 0.0142f
C9301 VDD.t190 VSUBS 0.0114f
C9302 VDD.t346 VSUBS 0.0114f
C9303 VDD.n2169 VSUBS 0.0268f
C9304 VDD.n2170 VSUBS 0.0129f
C9305 VDD.n2171 VSUBS 0.00717f
C9306 VDD.n2172 VSUBS 0.00349f
C9307 VDD.n2173 VSUBS 0.0145f
C9308 VDD.n2174 VSUBS 0.0273f
C9309 VDD.n2175 VSUBS 0.0142f
C9310 VDD.t345 VSUBS 0.0114f
C9311 VDD.t227 VSUBS 0.0114f
C9312 VDD.n2176 VSUBS 0.0268f
C9313 VDD.n2177 VSUBS 0.0129f
C9314 VDD.n2178 VSUBS 0.00717f
C9315 VDD.n2179 VSUBS 0.00349f
C9316 VDD.n2180 VSUBS 0.0145f
C9317 VDD.n2181 VSUBS 0.0273f
C9318 VDD.n2182 VSUBS 0.0142f
C9319 VDD.t272 VSUBS 0.0114f
C9320 VDD.t233 VSUBS 0.0114f
C9321 VDD.n2183 VSUBS 0.0268f
C9322 VDD.n2184 VSUBS 0.0129f
C9323 VDD.n2185 VSUBS 0.00717f
C9324 VDD.n2186 VSUBS 0.00349f
C9325 VDD.n2187 VSUBS 0.0145f
C9326 VDD.n2188 VSUBS 0.0273f
C9327 VDD.n2189 VSUBS 0.0142f
C9328 VDD.t171 VSUBS 0.0114f
C9329 VDD.t321 VSUBS 0.0114f
C9330 VDD.n2190 VSUBS 0.0268f
C9331 VDD.n2191 VSUBS 0.0129f
C9332 VDD.n2192 VSUBS 0.00717f
C9333 VDD.n2193 VSUBS 0.00349f
C9334 VDD.n2194 VSUBS 0.0145f
C9335 VDD.n2195 VSUBS 0.0273f
C9336 VDD.n2196 VSUBS 0.0142f
C9337 VDD.t179 VSUBS 0.0114f
C9338 VDD.t217 VSUBS 0.0114f
C9339 VDD.n2197 VSUBS 0.0268f
C9340 VDD.n2198 VSUBS 0.0129f
C9341 VDD.n2199 VSUBS 0.00717f
C9342 VDD.n2200 VSUBS 0.00349f
C9343 VDD.n2201 VSUBS 0.0145f
C9344 VDD.n2202 VSUBS 0.0273f
C9345 VDD.n2203 VSUBS 0.0142f
C9346 VDD.t312 VSUBS 0.0114f
C9347 VDD.t222 VSUBS 0.0114f
C9348 VDD.n2204 VSUBS 0.0268f
C9349 VDD.n2205 VSUBS 0.0129f
C9350 VDD.n2206 VSUBS 0.00717f
C9351 VDD.n2207 VSUBS 0.00349f
C9352 VDD.n2208 VSUBS 0.0145f
C9353 VDD.n2209 VSUBS 0.0273f
C9354 VDD.n2210 VSUBS 0.0142f
C9355 VDD.t356 VSUBS 0.0114f
C9356 VDD.t305 VSUBS 0.0114f
C9357 VDD.n2211 VSUBS 0.0268f
C9358 VDD.n2212 VSUBS 0.0129f
C9359 VDD.n2213 VSUBS 0.00717f
C9360 VDD.n2214 VSUBS 0.00349f
C9361 VDD.n2215 VSUBS 0.0145f
C9362 VDD.n2216 VSUBS 0.0273f
C9363 VDD.n2217 VSUBS 0.0142f
C9364 VDD.t295 VSUBS 0.0114f
C9365 VDD.t241 VSUBS 0.0114f
C9366 VDD.n2218 VSUBS 0.0268f
C9367 VDD.n2219 VSUBS 0.0129f
C9368 VDD.n2220 VSUBS 0.00717f
C9369 VDD.n2221 VSUBS 0.00349f
C9370 VDD.n2222 VSUBS 0.0145f
C9371 VDD.n2223 VSUBS 0.0273f
C9372 VDD.n2224 VSUBS 0.0142f
C9373 VDD.t193 VSUBS 0.0114f
C9374 VDD.t201 VSUBS 0.0114f
C9375 VDD.n2225 VSUBS 0.0268f
C9376 VDD.n2226 VSUBS 0.0129f
C9377 VDD.n2227 VSUBS 0.00717f
C9378 VDD.n2228 VSUBS 0.00349f
C9379 VDD.n2229 VSUBS 0.0145f
C9380 VDD.n2230 VSUBS 0.0273f
C9381 VDD.n2231 VSUBS 0.0142f
C9382 VDD.t328 VSUBS 0.0114f
C9383 VDD.t276 VSUBS 0.0114f
C9384 VDD.n2232 VSUBS 0.0268f
C9385 VDD.n2233 VSUBS 0.0129f
C9386 VDD.n2234 VSUBS 0.00717f
C9387 VDD.n2235 VSUBS 0.00349f
C9388 VDD.n2236 VSUBS 0.0145f
C9389 VDD.n2237 VSUBS 0.0273f
C9390 VDD.n2238 VSUBS 0.0142f
C9391 VDD.t300 VSUBS 0.0114f
C9392 VDD.t176 VSUBS 0.0114f
C9393 VDD.n2239 VSUBS 0.0268f
C9394 VDD.n2240 VSUBS 0.0129f
C9395 VDD.n2241 VSUBS 0.00717f
C9396 VDD.n2242 VSUBS 0.00349f
C9397 VDD.n2243 VSUBS 0.0145f
C9398 VDD.n2244 VSUBS 0.0273f
C9399 VDD.n2245 VSUBS 0.0142f
C9400 VDD.t357 VSUBS 0.0114f
C9401 VDD.t242 VSUBS 0.0114f
C9402 VDD.n2246 VSUBS 0.0268f
C9403 VDD.n2247 VSUBS 0.0129f
C9404 VDD.n2248 VSUBS 0.00717f
C9405 VDD.n2249 VSUBS 0.00349f
C9406 VDD.n2250 VSUBS 0.0145f
C9407 VDD.n2251 VSUBS 0.0273f
C9408 VDD.n2252 VSUBS 0.0142f
C9409 VDD.t256 VSUBS 0.0114f
C9410 VDD.t307 VSUBS 0.0114f
C9411 VDD.n2253 VSUBS 0.0268f
C9412 VDD.n2254 VSUBS 0.0129f
C9413 VDD.n2255 VSUBS 0.00717f
C9414 VDD.n2256 VSUBS 0.00349f
C9415 VDD.n2257 VSUBS 0.0145f
C9416 VDD.n2258 VSUBS 0.0273f
C9417 VDD.n2259 VSUBS 0.0142f
C9418 VDD.t180 VSUBS 0.0114f
C9419 VDD.t172 VSUBS 0.0114f
C9420 VDD.n2260 VSUBS 0.0268f
C9421 VDD.n2261 VSUBS 0.0129f
C9422 VDD.n2262 VSUBS 0.00717f
C9423 VDD.n2263 VSUBS 0.00349f
C9424 VDD.n2264 VSUBS 0.0145f
C9425 VDD.n2265 VSUBS 0.0273f
C9426 VDD.n2266 VSUBS 0.0142f
C9427 VDD.t239 VSUBS 0.0114f
C9428 VDD.t279 VSUBS 0.0114f
C9429 VDD.n2267 VSUBS 0.0268f
C9430 VDD.n2268 VSUBS 0.0129f
C9431 VDD.n2269 VSUBS 0.00717f
C9432 VDD.n2270 VSUBS 0.00349f
C9433 VDD.n2271 VSUBS 0.0145f
C9434 VDD.n2272 VSUBS 0.0273f
C9435 VDD.n2273 VSUBS 0.0142f
C9436 VDD.t296 VSUBS 0.0114f
C9437 VDD.t350 VSUBS 0.0114f
C9438 VDD.n2274 VSUBS 0.0268f
C9439 VDD.n2275 VSUBS 0.0129f
C9440 VDD.n2276 VSUBS 0.00717f
C9441 VDD.n2277 VSUBS 0.00349f
C9442 VDD.n2278 VSUBS 0.0145f
C9443 VDD.n2279 VSUBS 0.0273f
C9444 VDD.n2280 VSUBS 0.0142f
C9445 VDD.t219 VSUBS 0.0114f
C9446 VDD.t309 VSUBS 0.0114f
C9447 VDD.n2281 VSUBS 0.0268f
C9448 VDD.n2282 VSUBS 0.0129f
C9449 VDD.n2283 VSUBS 0.00717f
C9450 VDD.n2284 VSUBS 0.00349f
C9451 VDD.n2285 VSUBS 0.0145f
C9452 VDD.n2286 VSUBS 0.0273f
C9453 VDD.n2287 VSUBS 0.0142f
C9454 VDD.t212 VSUBS 0.0114f
C9455 VDD.t299 VSUBS 0.0114f
C9456 VDD.n2288 VSUBS 0.0268f
C9457 VDD.n2289 VSUBS 0.0129f
C9458 VDD.n2290 VSUBS 0.00717f
C9459 VDD.n2291 VSUBS 0.00349f
C9460 VDD.n2292 VSUBS 0.0202f
C9461 VDD.n2293 VSUBS 0.0273f
C9462 VDD.n2294 VSUBS 0.0142f
C9463 VDD.n2295 VSUBS 0.215f
C9464 VDD.n2296 VSUBS 0.0867f
C9465 VDD.n2297 VSUBS 0.0867f
C9466 VDD.n2298 VSUBS 0.0867f
C9467 VDD.n2299 VSUBS 0.0867f
C9468 VDD.n2300 VSUBS 0.0867f
C9469 VDD.n2301 VSUBS 0.0867f
C9470 VDD.n2302 VSUBS 0.0867f
C9471 VDD.n2303 VSUBS 0.0867f
C9472 VDD.n2304 VSUBS 0.0867f
C9473 VDD.n2305 VSUBS 0.0867f
C9474 VDD.n2306 VSUBS 0.0867f
C9475 VDD.n2307 VSUBS 0.0867f
C9476 VDD.n2308 VSUBS 0.0867f
C9477 VDD.n2309 VSUBS 0.0867f
C9478 VDD.n2310 VSUBS 0.0867f
C9479 VDD.n2311 VSUBS 0.0867f
C9480 VDD.n2312 VSUBS 0.0867f
C9481 VDD.n2313 VSUBS 0.0867f
C9482 VDD.n2314 VSUBS 0.0867f
C9483 VDD.n2315 VSUBS 0.0867f
C9484 VDD.n2316 VSUBS 0.0867f
C9485 VDD.n2317 VSUBS 0.0867f
C9486 VDD.n2318 VSUBS 0.0867f
C9487 VDD.n2319 VSUBS 0.0867f
C9488 VDD.n2320 VSUBS 0.0867f
C9489 VDD.n2321 VSUBS 0.0867f
C9490 VDD.n2322 VSUBS 0.0867f
C9491 VDD.n2323 VSUBS 0.0867f
C9492 VDD.n2324 VSUBS 0.0867f
C9493 VDD.n2325 VSUBS 0.0867f
C9494 VDD.n2326 VSUBS 0.0867f
C9495 VDD.n2327 VSUBS 0.0867f
C9496 VDD.n2328 VSUBS 0.0867f
C9497 VDD.n2329 VSUBS 0.0867f
C9498 VDD.n2330 VSUBS 0.0867f
C9499 VDD.n2331 VSUBS 0.0867f
C9500 VDD.n2332 VSUBS 0.0867f
C9501 VDD.n2333 VSUBS 0.0867f
C9502 VDD.t310 VSUBS 0.0114f
C9503 VDD.t261 VSUBS 0.0114f
C9504 VDD.n2334 VSUBS 0.0269f
C9505 VDD.n2335 VSUBS 0.0132f
C9506 VDD.n2336 VSUBS 0.0071f
C9507 VDD.n2337 VSUBS 0.00345f
C9508 VDD.n2338 VSUBS 0.0145f
C9509 VDD.n2339 VSUBS 0.0275f
C9510 VDD.n2340 VSUBS 0.0142f
C9511 VDD.t244 VSUBS 0.0114f
C9512 VDD.t361 VSUBS 0.0114f
C9513 VDD.n2341 VSUBS 0.0269f
C9514 VDD.n2342 VSUBS 0.0132f
C9515 VDD.n2343 VSUBS 0.0071f
C9516 VDD.n2344 VSUBS 0.00345f
C9517 VDD.n2345 VSUBS 0.0145f
C9518 VDD.n2346 VSUBS 0.0275f
C9519 VDD.n2347 VSUBS 0.0142f
C9520 VDD.t342 VSUBS 0.0114f
C9521 VDD.t290 VSUBS 0.0114f
C9522 VDD.n2348 VSUBS 0.0269f
C9523 VDD.n2349 VSUBS 0.0132f
C9524 VDD.n2350 VSUBS 0.0071f
C9525 VDD.n2351 VSUBS 0.00345f
C9526 VDD.n2352 VSUBS 0.0145f
C9527 VDD.n2353 VSUBS 0.0275f
C9528 VDD.n2354 VSUBS 0.0142f
C9529 VDD.t288 VSUBS 0.0114f
C9530 VDD.t188 VSUBS 0.0114f
C9531 VDD.n2355 VSUBS 0.0269f
C9532 VDD.n2356 VSUBS 0.0132f
C9533 VDD.n2357 VSUBS 0.0071f
C9534 VDD.n2358 VSUBS 0.00345f
C9535 VDD.n2359 VSUBS 0.0145f
C9536 VDD.n2360 VSUBS 0.0275f
C9537 VDD.n2361 VSUBS 0.0142f
C9538 VDD.t232 VSUBS 0.0114f
C9539 VDD.t195 VSUBS 0.0114f
C9540 VDD.n2362 VSUBS 0.0269f
C9541 VDD.n2363 VSUBS 0.0132f
C9542 VDD.n2364 VSUBS 0.0071f
C9543 VDD.n2365 VSUBS 0.00345f
C9544 VDD.n2366 VSUBS 0.0145f
C9545 VDD.n2367 VSUBS 0.0275f
C9546 VDD.n2368 VSUBS 0.0142f
C9547 VDD.t318 VSUBS 0.0114f
C9548 VDD.t271 VSUBS 0.0114f
C9549 VDD.n2369 VSUBS 0.0269f
C9550 VDD.n2370 VSUBS 0.0132f
C9551 VDD.n2371 VSUBS 0.0071f
C9552 VDD.n2372 VSUBS 0.00345f
C9553 VDD.n2373 VSUBS 0.0145f
C9554 VDD.n2374 VSUBS 0.0275f
C9555 VDD.n2375 VSUBS 0.0142f
C9556 VDD.t330 VSUBS 0.0114f
C9557 VDD.t168 VSUBS 0.0114f
C9558 VDD.n2376 VSUBS 0.0269f
C9559 VDD.n2377 VSUBS 0.0132f
C9560 VDD.n2378 VSUBS 0.0071f
C9561 VDD.n2379 VSUBS 0.00345f
C9562 VDD.n2380 VSUBS 0.0145f
C9563 VDD.n2381 VSUBS 0.0275f
C9564 VDD.n2382 VSUBS 0.0142f
C9565 VDD.t259 VSUBS 0.0114f
C9566 VDD.t177 VSUBS 0.0114f
C9567 VDD.n2383 VSUBS 0.0269f
C9568 VDD.n2384 VSUBS 0.0132f
C9569 VDD.n2385 VSUBS 0.0071f
C9570 VDD.n2386 VSUBS 0.00345f
C9571 VDD.n2387 VSUBS 0.0145f
C9572 VDD.n2388 VSUBS 0.0275f
C9573 VDD.n2389 VSUBS 0.0142f
C9574 VDD.t302 VSUBS 0.0114f
C9575 VDD.t254 VSUBS 0.0114f
C9576 VDD.n2390 VSUBS 0.0269f
C9577 VDD.n2391 VSUBS 0.0132f
C9578 VDD.n2392 VSUBS 0.0071f
C9579 VDD.n2393 VSUBS 0.00345f
C9580 VDD.n2394 VSUBS 0.0145f
C9581 VDD.n2395 VSUBS 0.0275f
C9582 VDD.n2396 VSUBS 0.0142f
C9583 VDD.t247 VSUBS 0.0114f
C9584 VDD.t203 VSUBS 0.0114f
C9585 VDD.n2397 VSUBS 0.0269f
C9586 VDD.n2398 VSUBS 0.0132f
C9587 VDD.n2399 VSUBS 0.0071f
C9588 VDD.n2400 VSUBS 0.00345f
C9589 VDD.n2401 VSUBS 0.0145f
C9590 VDD.n2402 VSUBS 0.0275f
C9591 VDD.n2403 VSUBS 0.0142f
C9592 VDD.t344 VSUBS 0.0114f
C9593 VDD.t355 VSUBS 0.0114f
C9594 VDD.n2404 VSUBS 0.0269f
C9595 VDD.n2405 VSUBS 0.0132f
C9596 VDD.n2406 VSUBS 0.0071f
C9597 VDD.n2407 VSUBS 0.00345f
C9598 VDD.n2408 VSUBS 0.0145f
C9599 VDD.n2409 VSUBS 0.0275f
C9600 VDD.n2410 VSUBS 0.0142f
C9601 VDD.t275 VSUBS 0.0114f
C9602 VDD.t236 VSUBS 0.0114f
C9603 VDD.n2411 VSUBS 0.0269f
C9604 VDD.n2412 VSUBS 0.0132f
C9605 VDD.n2413 VSUBS 0.0071f
C9606 VDD.n2414 VSUBS 0.00345f
C9607 VDD.n2415 VSUBS 0.0145f
C9608 VDD.n2416 VSUBS 0.0275f
C9609 VDD.n2417 VSUBS 0.0142f
C9610 VDD.t251 VSUBS 0.0114f
C9611 VDD.t324 VSUBS 0.0114f
C9612 VDD.n2418 VSUBS 0.0269f
C9613 VDD.n2419 VSUBS 0.0132f
C9614 VDD.n2420 VSUBS 0.0071f
C9615 VDD.n2421 VSUBS 0.00345f
C9616 VDD.n2422 VSUBS 0.0145f
C9617 VDD.n2423 VSUBS 0.0275f
C9618 VDD.n2424 VSUBS 0.0142f
C9619 VDD.t303 VSUBS 0.0114f
C9620 VDD.t205 VSUBS 0.0114f
C9621 VDD.n2425 VSUBS 0.0269f
C9622 VDD.n2426 VSUBS 0.0132f
C9623 VDD.n2427 VSUBS 0.0071f
C9624 VDD.n2428 VSUBS 0.00345f
C9625 VDD.n2429 VSUBS 0.0145f
C9626 VDD.n2430 VSUBS 0.0275f
C9627 VDD.n2431 VSUBS 0.0142f
C9628 VDD.t221 VSUBS 0.0114f
C9629 VDD.t250 VSUBS 0.0114f
C9630 VDD.n2432 VSUBS 0.0269f
C9631 VDD.n2433 VSUBS 0.0132f
C9632 VDD.n2434 VSUBS 0.0071f
C9633 VDD.n2435 VSUBS 0.00345f
C9634 VDD.n2436 VSUBS 0.0145f
C9635 VDD.n2437 VSUBS 0.0275f
C9636 VDD.n2438 VSUBS 0.0142f
C9637 VDD.t331 VSUBS 0.0114f
C9638 VDD.t319 VSUBS 0.0114f
C9639 VDD.n2439 VSUBS 0.0269f
C9640 VDD.n2440 VSUBS 0.0132f
C9641 VDD.n2441 VSUBS 0.0071f
C9642 VDD.n2442 VSUBS 0.00345f
C9643 VDD.n2443 VSUBS 0.0145f
C9644 VDD.n2444 VSUBS 0.0275f
C9645 VDD.n2445 VSUBS 0.0142f
C9646 VDD.t199 VSUBS 0.0114f
C9647 VDD.t237 VSUBS 0.0114f
C9648 VDD.n2446 VSUBS 0.0269f
C9649 VDD.n2447 VSUBS 0.0132f
C9650 VDD.n2448 VSUBS 0.0071f
C9651 VDD.n2449 VSUBS 0.00345f
C9652 VDD.n2450 VSUBS 0.0145f
C9653 VDD.n2451 VSUBS 0.0275f
C9654 VDD.n2452 VSUBS 0.0142f
C9655 VDD.t248 VSUBS 0.0114f
C9656 VDD.t294 VSUBS 0.0114f
C9657 VDD.n2453 VSUBS 0.0269f
C9658 VDD.n2454 VSUBS 0.0132f
C9659 VDD.n2455 VSUBS 0.0071f
C9660 VDD.n2456 VSUBS 0.00345f
C9661 VDD.n2457 VSUBS 0.0145f
C9662 VDD.n2458 VSUBS 0.0275f
C9663 VDD.n2459 VSUBS 0.0142f
C9664 VDD.t173 VSUBS 0.0114f
C9665 VDD.t257 VSUBS 0.0114f
C9666 VDD.n2460 VSUBS 0.0269f
C9667 VDD.n2461 VSUBS 0.0132f
C9668 VDD.n2462 VSUBS 0.0071f
C9669 VDD.n2463 VSUBS 0.00345f
C9670 VDD.n2464 VSUBS 0.0145f
C9671 VDD.n2465 VSUBS 0.0275f
C9672 VDD.n2466 VSUBS 0.0142f
C9673 VDD.t365 VSUBS 0.0114f
C9674 VDD.t249 VSUBS 0.0114f
C9675 VDD.n2467 VSUBS 0.0269f
C9676 VDD.n2468 VSUBS 0.0132f
C9677 VDD.n2469 VSUBS 0.0071f
C9678 VDD.n2470 VSUBS 0.00345f
C9679 VDD.n2471 VSUBS 0.0202f
C9680 VDD.n2472 VSUBS 0.0275f
C9681 VDD.n2473 VSUBS 0.0142f
C9682 VDD.n2474 VSUBS 0.215f
C9683 VDD.n2475 VSUBS 0.0867f
C9684 VDD.n2476 VSUBS 0.0867f
C9685 VDD.n2477 VSUBS 0.0867f
C9686 VDD.n2478 VSUBS 0.0867f
C9687 VDD.n2479 VSUBS 0.0867f
C9688 VDD.n2480 VSUBS 0.0867f
C9689 VDD.n2481 VSUBS 0.0867f
C9690 VDD.n2482 VSUBS 0.0867f
C9691 VDD.n2483 VSUBS 0.0867f
C9692 VDD.n2484 VSUBS 0.0867f
C9693 VDD.n2485 VSUBS 0.0867f
C9694 VDD.n2486 VSUBS 0.0867f
C9695 VDD.n2487 VSUBS 0.0867f
C9696 VDD.n2488 VSUBS 0.0867f
C9697 VDD.n2489 VSUBS 0.0867f
C9698 VDD.n2490 VSUBS 0.0867f
C9699 VDD.n2491 VSUBS 0.0867f
C9700 VDD.n2492 VSUBS 0.0867f
C9701 VDD.n2493 VSUBS 0.0867f
C9702 VDD.n2494 VSUBS 0.0867f
C9703 VDD.n2495 VSUBS 0.0867f
C9704 VDD.n2496 VSUBS 0.0867f
C9705 VDD.n2497 VSUBS 0.0867f
C9706 VDD.n2498 VSUBS 0.0867f
C9707 VDD.n2499 VSUBS 0.0867f
C9708 VDD.n2500 VSUBS 0.0867f
C9709 VDD.n2501 VSUBS 0.0867f
C9710 VDD.n2502 VSUBS 0.0867f
C9711 VDD.n2503 VSUBS 0.0867f
C9712 VDD.n2504 VSUBS 0.0867f
C9713 VDD.n2505 VSUBS 0.0867f
C9714 VDD.n2506 VSUBS 0.0867f
C9715 VDD.n2507 VSUBS 0.0867f
C9716 VDD.n2508 VSUBS 0.0867f
C9717 VDD.n2509 VSUBS 0.0867f
C9718 VDD.n2510 VSUBS 0.0867f
C9719 VDD.n2511 VSUBS 0.0867f
C9720 VDD.n2512 VSUBS 0.0867f
C9721 VDD.t186 VSUBS 0.0114f
C9722 VDD.t343 VSUBS 0.0114f
C9723 VDD.n2513 VSUBS 0.0269f
C9724 VDD.n2514 VSUBS 0.0133f
C9725 VDD.n2515 VSUBS 0.0071f
C9726 VDD.n2516 VSUBS 0.00345f
C9727 VDD.n2517 VSUBS 0.0145f
C9728 VDD.n2518 VSUBS 0.0275f
C9729 VDD.n2519 VSUBS 0.0142f
C9730 VDD.t320 VSUBS 0.0114f
C9731 VDD.t226 VSUBS 0.0114f
C9732 VDD.n2520 VSUBS 0.0269f
C9733 VDD.n2521 VSUBS 0.0133f
C9734 VDD.n2522 VSUBS 0.0071f
C9735 VDD.n2523 VSUBS 0.00345f
C9736 VDD.n2524 VSUBS 0.0145f
C9737 VDD.n2525 VSUBS 0.0275f
C9738 VDD.n2526 VSUBS 0.0142f
C9739 VDD.t214 VSUBS 0.0114f
C9740 VDD.t170 VSUBS 0.0114f
C9741 VDD.n2527 VSUBS 0.0269f
C9742 VDD.n2528 VSUBS 0.0133f
C9743 VDD.n2529 VSUBS 0.0071f
C9744 VDD.n2530 VSUBS 0.00345f
C9745 VDD.n2531 VSUBS 0.0145f
C9746 VDD.n2532 VSUBS 0.0275f
C9747 VDD.n2533 VSUBS 0.0142f
C9748 VDD.t169 VSUBS 0.0114f
C9749 VDD.t245 VSUBS 0.0114f
C9750 VDD.n2534 VSUBS 0.0269f
C9751 VDD.n2535 VSUBS 0.0133f
C9752 VDD.n2536 VSUBS 0.0071f
C9753 VDD.n2537 VSUBS 0.00345f
C9754 VDD.n2538 VSUBS 0.0145f
C9755 VDD.n2539 VSUBS 0.0275f
C9756 VDD.n2540 VSUBS 0.0142f
C9757 VDD.t304 VSUBS 0.0114f
C9758 VDD.t255 VSUBS 0.0114f
C9759 VDD.n2541 VSUBS 0.0269f
C9760 VDD.n2542 VSUBS 0.0133f
C9761 VDD.n2543 VSUBS 0.0071f
C9762 VDD.n2544 VSUBS 0.00345f
C9763 VDD.n2545 VSUBS 0.0145f
C9764 VDD.n2546 VSUBS 0.0275f
C9765 VDD.n2547 VSUBS 0.0142f
C9766 VDD.t191 VSUBS 0.0114f
C9767 VDD.t354 VSUBS 0.0114f
C9768 VDD.n2548 VSUBS 0.0269f
C9769 VDD.n2549 VSUBS 0.0133f
C9770 VDD.n2550 VSUBS 0.0071f
C9771 VDD.n2551 VSUBS 0.00345f
C9772 VDD.n2552 VSUBS 0.0145f
C9773 VDD.n2553 VSUBS 0.0275f
C9774 VDD.n2554 VSUBS 0.0142f
C9775 VDD.t204 VSUBS 0.0114f
C9776 VDD.t235 VSUBS 0.0114f
C9777 VDD.n2555 VSUBS 0.0269f
C9778 VDD.n2556 VSUBS 0.0133f
C9779 VDD.n2557 VSUBS 0.0071f
C9780 VDD.n2558 VSUBS 0.00345f
C9781 VDD.n2559 VSUBS 0.0145f
C9782 VDD.n2560 VSUBS 0.0275f
C9783 VDD.n2561 VSUBS 0.0142f
C9784 VDD.t340 VSUBS 0.0114f
C9785 VDD.t240 VSUBS 0.0114f
C9786 VDD.n2562 VSUBS 0.0269f
C9787 VDD.n2563 VSUBS 0.0133f
C9788 VDD.n2564 VSUBS 0.0071f
C9789 VDD.n2565 VSUBS 0.00345f
C9790 VDD.n2566 VSUBS 0.0145f
C9791 VDD.n2567 VSUBS 0.0275f
C9792 VDD.n2568 VSUBS 0.0142f
C9793 VDD.t182 VSUBS 0.0114f
C9794 VDD.t334 VSUBS 0.0114f
C9795 VDD.n2569 VSUBS 0.0269f
C9796 VDD.n2570 VSUBS 0.0133f
C9797 VDD.n2571 VSUBS 0.0071f
C9798 VDD.n2572 VSUBS 0.00345f
C9799 VDD.n2573 VSUBS 0.0145f
C9800 VDD.n2574 VSUBS 0.0275f
C9801 VDD.n2575 VSUBS 0.0142f
C9802 VDD.t325 VSUBS 0.0114f
C9803 VDD.t262 VSUBS 0.0114f
C9804 VDD.n2576 VSUBS 0.0269f
C9805 VDD.n2577 VSUBS 0.0133f
C9806 VDD.n2578 VSUBS 0.0071f
C9807 VDD.n2579 VSUBS 0.00345f
C9808 VDD.n2580 VSUBS 0.0145f
C9809 VDD.n2581 VSUBS 0.0275f
C9810 VDD.n2582 VSUBS 0.0142f
C9811 VDD.t218 VSUBS 0.0114f
C9812 VDD.t216 VSUBS 0.0114f
C9813 VDD.n2583 VSUBS 0.0269f
C9814 VDD.n2584 VSUBS 0.0133f
C9815 VDD.n2585 VSUBS 0.0071f
C9816 VDD.n2586 VSUBS 0.00345f
C9817 VDD.n2587 VSUBS 0.0145f
C9818 VDD.n2588 VSUBS 0.0275f
C9819 VDD.n2589 VSUBS 0.0142f
C9820 VDD.t358 VSUBS 0.0114f
C9821 VDD.t308 VSUBS 0.0114f
C9822 VDD.n2590 VSUBS 0.0269f
C9823 VDD.n2591 VSUBS 0.0133f
C9824 VDD.n2592 VSUBS 0.0071f
C9825 VDD.n2593 VSUBS 0.00345f
C9826 VDD.n2594 VSUBS 0.0145f
C9827 VDD.n2595 VSUBS 0.0275f
C9828 VDD.n2596 VSUBS 0.0142f
C9829 VDD.t329 VSUBS 0.0114f
C9830 VDD.t202 VSUBS 0.0114f
C9831 VDD.n2597 VSUBS 0.0269f
C9832 VDD.n2598 VSUBS 0.0133f
C9833 VDD.n2599 VSUBS 0.0071f
C9834 VDD.n2600 VSUBS 0.00345f
C9835 VDD.n2601 VSUBS 0.0145f
C9836 VDD.n2602 VSUBS 0.0275f
C9837 VDD.n2603 VSUBS 0.0142f
C9838 VDD.t184 VSUBS 0.0114f
C9839 VDD.t263 VSUBS 0.0114f
C9840 VDD.n2604 VSUBS 0.0269f
C9841 VDD.n2605 VSUBS 0.0133f
C9842 VDD.n2606 VSUBS 0.0071f
C9843 VDD.n2607 VSUBS 0.00345f
C9844 VDD.n2608 VSUBS 0.0145f
C9845 VDD.n2609 VSUBS 0.0275f
C9846 VDD.n2610 VSUBS 0.0142f
C9847 VDD.t280 VSUBS 0.0114f
C9848 VDD.t335 VSUBS 0.0114f
C9849 VDD.n2611 VSUBS 0.0269f
C9850 VDD.n2612 VSUBS 0.0133f
C9851 VDD.n2613 VSUBS 0.0071f
C9852 VDD.n2614 VSUBS 0.00345f
C9853 VDD.n2615 VSUBS 0.0145f
C9854 VDD.n2616 VSUBS 0.0275f
C9855 VDD.n2617 VSUBS 0.0142f
C9856 VDD.t207 VSUBS 0.0114f
C9857 VDD.t197 VSUBS 0.0114f
C9858 VDD.n2618 VSUBS 0.0269f
C9859 VDD.n2619 VSUBS 0.0133f
C9860 VDD.n2620 VSUBS 0.0071f
C9861 VDD.n2621 VSUBS 0.00345f
C9862 VDD.n2622 VSUBS 0.0145f
C9863 VDD.n2623 VSUBS 0.0275f
C9864 VDD.n2624 VSUBS 0.0142f
C9865 VDD.t258 VSUBS 0.0114f
C9866 VDD.t306 VSUBS 0.0114f
C9867 VDD.n2625 VSUBS 0.0269f
C9868 VDD.n2626 VSUBS 0.0133f
C9869 VDD.n2627 VSUBS 0.0071f
C9870 VDD.n2628 VSUBS 0.00345f
C9871 VDD.n2629 VSUBS 0.0145f
C9872 VDD.n2630 VSUBS 0.0275f
C9873 VDD.n2631 VSUBS 0.0142f
C9874 VDD.t326 VSUBS 0.0114f
C9875 VDD.t175 VSUBS 0.0114f
C9876 VDD.n2632 VSUBS 0.0269f
C9877 VDD.n2633 VSUBS 0.0133f
C9878 VDD.n2634 VSUBS 0.0071f
C9879 VDD.n2635 VSUBS 0.00345f
C9880 VDD.n2636 VSUBS 0.0145f
C9881 VDD.n2637 VSUBS 0.0275f
C9882 VDD.n2638 VSUBS 0.0142f
C9883 VDD.t238 VSUBS 0.0114f
C9884 VDD.t337 VSUBS 0.0114f
C9885 VDD.n2639 VSUBS 0.0269f
C9886 VDD.n2640 VSUBS 0.0133f
C9887 VDD.n2641 VSUBS 0.0071f
C9888 VDD.n2642 VSUBS 0.00345f
C9889 VDD.n2643 VSUBS 0.0145f
C9890 VDD.n2644 VSUBS 0.0275f
C9891 VDD.n2645 VSUBS 0.0142f
C9892 VDD.t229 VSUBS 0.0114f
C9893 VDD.t327 VSUBS 0.0114f
C9894 VDD.n2646 VSUBS 0.0269f
C9895 VDD.n2647 VSUBS 0.0133f
C9896 VDD.n2648 VSUBS 0.0071f
C9897 VDD.n2649 VSUBS 0.00345f
C9898 VDD.n2650 VSUBS 0.0202f
C9899 VDD.n2651 VSUBS 0.0275f
C9900 VDD.n2652 VSUBS 0.0142f
C9901 VDD.n2653 VSUBS 0.215f
C9902 VDD.n2654 VSUBS 0.0867f
C9903 VDD.n2655 VSUBS 0.0867f
C9904 VDD.n2656 VSUBS 0.0867f
C9905 VDD.n2657 VSUBS 0.0867f
C9906 VDD.n2658 VSUBS 0.0867f
C9907 VDD.n2659 VSUBS 0.0867f
C9908 VDD.n2660 VSUBS 0.0867f
C9909 VDD.n2661 VSUBS 0.0867f
C9910 VDD.n2662 VSUBS 0.0867f
C9911 VDD.n2663 VSUBS 0.0867f
C9912 VDD.n2664 VSUBS 0.0867f
C9913 VDD.n2665 VSUBS 0.0867f
C9914 VDD.n2666 VSUBS 0.0867f
C9915 VDD.n2667 VSUBS 0.0867f
C9916 VDD.n2668 VSUBS 0.0867f
C9917 VDD.n2669 VSUBS 0.0867f
C9918 VDD.n2670 VSUBS 0.0867f
C9919 VDD.n2671 VSUBS 0.0867f
C9920 VDD.n2672 VSUBS 0.0867f
C9921 VDD.n2673 VSUBS 0.0867f
C9922 VDD.n2674 VSUBS 0.0867f
C9923 VDD.n2675 VSUBS 0.0867f
C9924 VDD.n2676 VSUBS 0.0867f
C9925 VDD.n2677 VSUBS 0.0867f
C9926 VDD.n2678 VSUBS 0.0867f
C9927 VDD.n2679 VSUBS 0.0867f
C9928 VDD.n2680 VSUBS 0.0867f
C9929 VDD.n2681 VSUBS 0.0867f
C9930 VDD.n2682 VSUBS 0.0867f
C9931 VDD.n2683 VSUBS 0.0867f
C9932 VDD.n2684 VSUBS 0.0867f
C9933 VDD.n2685 VSUBS 0.0867f
C9934 VDD.n2686 VSUBS 0.0867f
C9935 VDD.n2687 VSUBS 0.0867f
C9936 VDD.n2688 VSUBS 0.0867f
C9937 VDD.n2689 VSUBS 0.0867f
C9938 VDD.n2690 VSUBS 0.0867f
C9939 VDD.n2691 VSUBS 0.0867f
C9940 VDD.n2692 VSUBS 0.0198f
C9941 VDD.n2693 VSUBS 0.0688f
C9942 VDD.n2694 VSUBS 0.0836f
C9943 VDD.n2695 VSUBS 0.0421f
C9944 VDD.n2696 VSUBS 0.0421f
C9945 VDD.n2697 VSUBS 0.0533f
C9946 VDD.n2698 VSUBS 0.0842f
C9947 VDD.n2699 VSUBS 0.0842f
C9948 VDD.n2700 VSUBS 0.0483f
C9949 VDD.n2701 VSUBS 0.0671f
C9950 VDD.n2702 VSUBS 0.0614f
C9951 VDD.n2703 VSUBS 0.0405f
C9952 VDD.n2704 VSUBS 0.0405f
C9953 VDD.n2705 VSUBS 0.0405f
C9954 VDD.n2706 VSUBS 0.0405f
C9955 VDD.n2707 VSUBS 0.0405f
C9956 VDD.n2708 VSUBS 0.0405f
C9957 VDD.n2709 VSUBS 0.0405f
C9958 VDD.n2710 VSUBS 0.0405f
C9959 VDD.n2711 VSUBS 0.0405f
C9960 VDD.n2712 VSUBS 0.0405f
C9961 VDD.n2713 VSUBS 0.0405f
C9962 VDD.n2714 VSUBS 0.0405f
C9963 VDD.n2715 VSUBS 0.0405f
C9964 VDD.n2716 VSUBS 0.0405f
C9965 VDD.n2717 VSUBS 0.0405f
C9966 VDD.n2718 VSUBS 0.0405f
C9967 VDD.n2719 VSUBS 0.0405f
C9968 VDD.n2720 VSUBS 0.0405f
C9969 VDD.n2721 VSUBS 0.0405f
C9970 VDD.n2722 VSUBS 0.0405f
C9971 VDD.n2723 VSUBS 0.0405f
C9972 VDD.n2724 VSUBS 0.0405f
C9973 VDD.n2725 VSUBS 0.0405f
C9974 VDD.n2726 VSUBS 0.0405f
C9975 VDD.n2727 VSUBS 0.0405f
C9976 VDD.n2728 VSUBS 0.0405f
C9977 VDD.n2729 VSUBS 0.0405f
C9978 VDD.n2730 VSUBS 0.0405f
C9979 VDD.n2731 VSUBS 0.0405f
C9980 VDD.n2732 VSUBS 0.0198f
C9981 VDD.n2733 VSUBS 0.0405f
C9982 VDD.n2734 VSUBS 0.0405f
C9983 VDD.n2735 VSUBS 0.0198f
C9984 VDD.n2736 VSUBS 0.0405f
C9985 VDD.n2737 VSUBS 0.0405f
C9986 VDD.n2738 VSUBS 0.0198f
C9987 VDD.n2739 VSUBS 0.0405f
C9988 VDD.n2740 VSUBS 0.0405f
C9989 VDD.n2741 VSUBS 0.0198f
C9990 VDD.n2742 VSUBS 0.0405f
C9991 VDD.n2743 VSUBS 0.0405f
C9992 VDD.n2744 VSUBS 0.0198f
C9993 VDD.n2745 VSUBS 0.0405f
C9994 VDD.n2746 VSUBS 0.0405f
C9995 VDD.n2747 VSUBS 0.0198f
C9996 VDD.n2748 VSUBS 0.0405f
C9997 VDD.n2749 VSUBS 0.0405f
C9998 VDD.n2750 VSUBS 0.0198f
C9999 VDD.n2751 VSUBS 0.0405f
C10000 VDD.n2752 VSUBS 0.0405f
C10001 VDD.n2753 VSUBS 0.0198f
C10002 VDD.n2754 VSUBS 0.0405f
C10003 VDD.n2755 VSUBS 0.0405f
C10004 VDD.n2756 VSUBS 0.0198f
C10005 VDD.n2757 VSUBS 0.0405f
C10006 VDD.n2758 VSUBS 0.0405f
C10007 VDD.n2759 VSUBS 0.0198f
C10008 VDD.n2760 VSUBS 0.0405f
C10009 VDD.n2761 VSUBS 0.0405f
C10010 VDD.n2762 VSUBS 0.0198f
C10011 VDD.n2763 VSUBS 0.0405f
C10012 VDD.n2764 VSUBS 0.0405f
C10013 VDD.n2765 VSUBS 0.0198f
C10014 VDD.n2766 VSUBS 0.0405f
C10015 VDD.n2767 VSUBS 0.0405f
C10016 VDD.n2768 VSUBS 0.0198f
C10017 VDD.n2769 VSUBS 0.0405f
C10018 VDD.n2770 VSUBS 0.0405f
C10019 VDD.n2771 VSUBS 0.0198f
C10020 VDD.n2772 VSUBS 0.0405f
C10021 VDD.n2773 VSUBS 0.0405f
C10022 VDD.n2774 VSUBS 0.0198f
C10023 VDD.n2775 VSUBS 0.0405f
C10024 VDD.n2776 VSUBS 0.0405f
C10025 VDD.n2777 VSUBS 0.0198f
C10026 VDD.n2778 VSUBS 0.0405f
C10027 VDD.n2779 VSUBS 0.0405f
C10028 VDD.n2780 VSUBS 0.0198f
C10029 VDD.n2781 VSUBS 0.0405f
C10030 VDD.n2782 VSUBS 0.0181f
C10031 VDD.n2783 VSUBS 0.0405f
C10032 VDD.n2784 VSUBS 0.0198f
C10033 VDD.n2785 VSUBS 0.0447f
C10034 VDD.n2786 VSUBS 0.0198f
C10035 VDD.n2787 VSUBS 0.0673f
C10036 VDD.n2788 VSUBS 0.0405f
C10037 VDD.n2789 VSUBS 0.0198f
C10038 VDD.n2790 VSUBS 0.0405f
C10039 VDD.n2791 VSUBS 0.0405f
C10040 VDD.n2792 VSUBS 0.0198f
C10041 VDD.n2793 VSUBS 0.0405f
C10042 VDD.n2794 VSUBS 0.0405f
C10043 VDD.n2795 VSUBS 0.0198f
C10044 VDD.n2796 VSUBS 0.0405f
C10045 VDD.n2797 VSUBS 0.0405f
C10046 VDD.n2798 VSUBS 0.0198f
C10047 VDD.n2799 VSUBS 0.0405f
C10048 VDD.n2800 VSUBS 0.0405f
C10049 VDD.n2801 VSUBS 0.0198f
C10050 VDD.n2802 VSUBS 0.0405f
C10051 VDD.n2803 VSUBS 0.0405f
C10052 VDD.n2804 VSUBS 0.0198f
C10053 VDD.n2805 VSUBS 0.0405f
C10054 VDD.n2806 VSUBS 0.0405f
C10055 VDD.n2807 VSUBS 0.0198f
C10056 VDD.n2808 VSUBS 0.0405f
C10057 VDD.n2809 VSUBS 0.0405f
C10058 VDD.n2810 VSUBS 0.0198f
C10059 VDD.n2811 VSUBS 0.0405f
C10060 VDD.n2812 VSUBS 0.0405f
C10061 VDD.n2813 VSUBS 0.0198f
C10062 VDD.n2814 VSUBS 0.0405f
C10063 VDD.n2815 VSUBS 0.0405f
C10064 VDD.n2816 VSUBS 0.0198f
C10065 VDD.n2817 VSUBS 0.0405f
C10066 VDD.n2818 VSUBS 0.0405f
C10067 VDD.n2819 VSUBS 0.0198f
C10068 VDD.n2820 VSUBS 0.0405f
C10069 VDD.n2821 VSUBS 0.0405f
C10070 VDD.n2822 VSUBS 0.0198f
C10071 VDD.n2823 VSUBS 0.0405f
C10072 VDD.n2824 VSUBS 0.0405f
C10073 VDD.n2825 VSUBS 0.0198f
C10074 VDD.n2826 VSUBS 0.0405f
C10075 VDD.n2827 VSUBS 0.0181f
C10076 VDD.n2828 VSUBS 0.0405f
C10077 VDD.n2829 VSUBS 0.0198f
C10078 VDD.n2830 VSUBS 0.0578f
C10079 VDD.n2831 VSUBS 0.0198f
C10080 VDD.n2832 VSUBS 0.0542f
C10081 VDD.n2833 VSUBS 0.0449f
C10082 VDD.n2834 VSUBS 8.65e-19
C10083 VDD.n2835 VSUBS 0.0384f
C10084 VDD.n2836 VSUBS 0.00593f
C10085 VDD.n2837 VSUBS 0.00194f
C10086 VDD.n2838 VSUBS 0.0333f
C10087 VDD.n2839 VSUBS 0.00989f
C10088 VDD.n2840 VSUBS 0.0198f
C10089 VDD.n2841 VSUBS 0.00989f
C10090 VDD.n2868 VSUBS 0.0198f
C10091 VDD.n2870 VSUBS 0.0198f
C10092 VDD.n2871 VSUBS 0.0198f
C10093 VDD.n2873 VSUBS 0.0198f
C10094 VDD.n2874 VSUBS 0.0198f
C10095 VDD.n2876 VSUBS 0.0198f
C10096 VDD.n2877 VSUBS 0.0198f
C10097 VDD.n2879 VSUBS 0.0198f
C10098 VDD.n2880 VSUBS 0.0198f
C10099 VDD.n2882 VSUBS 0.0198f
C10100 VDD.n2883 VSUBS 0.0198f
C10101 VDD.n2885 VSUBS 0.0198f
C10102 VDD.n2886 VSUBS 0.0198f
C10103 VDD.n2888 VSUBS 0.0198f
C10104 VDD.n2889 VSUBS 0.0198f
C10105 VDD.n2891 VSUBS 2.66f
C10106 VDD.n2892 VSUBS 0.801f
C10107 VDD.n2893 VSUBS 0.0287f
C10108 VDD.n2894 VSUBS 0.916f
C10109 VDD.n2895 VSUBS 0.0198f
C10110 VDD.n2896 VSUBS 1.38f
C10111 VDD.n2897 VSUBS 0.0198f
C10112 VDD.n2898 VSUBS 1.26f
C10113 VDD.n2902 VSUBS 0.0155f
C10114 VDD.n2903 VSUBS 0.0155f
C10115 VDD.n2905 VSUBS 0.0155f
C10116 VDD.n2906 VSUBS 0.0155f
C10117 VDD.n2908 VSUBS 0.0155f
C10118 VDD.n2909 VSUBS 0.0155f
C10119 VDD.n2911 VSUBS 0.0155f
C10120 VDD.n2912 VSUBS 0.0155f
C10121 VDD.n2914 VSUBS 0.0155f
C10122 VDD.n2915 VSUBS 0.0155f
C10123 VDD.n2917 VSUBS 0.0155f
C10124 VDD.n2918 VSUBS 0.0155f
C10125 VDD.n2920 VSUBS 0.0155f
C10126 VDD.n2921 VSUBS 0.0155f
C10127 VDD.n2923 VSUBS 0.0155f
C10128 VDD.n2924 VSUBS 0.0155f
C10129 VDD.n2926 VSUBS 0.0155f
C10130 VDD.n2927 VSUBS 0.0155f
C10131 VDD.n2929 VSUBS 0.0155f
C10132 VDD.n2930 VSUBS 0.0155f
C10133 VDD.n2932 VSUBS 0.0155f
C10134 VDD.n2933 VSUBS 0.0155f
C10135 VDD.n2935 VSUBS 0.0155f
C10136 VDD.n2936 VSUBS 0.0155f
C10137 VDD.n2938 VSUBS 0.0155f
C10138 VDD.n2940 VSUBS 0.0155f
C10139 VDD.n2942 VSUBS 0.0155f
C10140 VDD.n2943 VSUBS 0.0155f
C10141 VDD.n2945 VSUBS 0.0155f
C10142 VDD.n2946 VSUBS 0.0155f
C10143 VDD.n2948 VSUBS 0.0155f
C10144 VDD.n2949 VSUBS 0.0155f
C10145 VDD.n2951 VSUBS 0.0155f
C10146 VDD.n2952 VSUBS 0.0155f
C10147 VDD.n2954 VSUBS 0.0155f
C10148 VDD.n2955 VSUBS 0.0155f
C10149 VDD.n2957 VSUBS 0.0155f
C10150 VDD.n2958 VSUBS 0.0155f
C10151 VDD.n2960 VSUBS 0.0155f
C10152 VDD.n2961 VSUBS 0.0155f
C10153 VDD.n2963 VSUBS 0.0155f
C10154 VDD.n2964 VSUBS 0.0155f
C10155 VDD.n2966 VSUBS 0.0155f
C10156 VDD.n2967 VSUBS 0.0155f
C10157 VDD.n2969 VSUBS 0.0155f
C10158 VDD.n2970 VSUBS 0.0155f
C10159 VDD.n2972 VSUBS 0.0155f
C10160 VDD.n2973 VSUBS 0.0155f
C10161 VDD.n2975 VSUBS 0.0155f
C10162 VDD.n2976 VSUBS 0.0155f
C10163 VDD.n2978 VSUBS 0.0155f
C10164 VDD.n2979 VSUBS 0.0155f
C10165 VDD.n2981 VSUBS 0.0155f
C10166 VDD.n2982 VSUBS 0.0155f
C10167 VDD.n2984 VSUBS 0.0155f
C10168 VDD.n2985 VSUBS 0.0327f
C10169 VDD.n2987 VSUBS 0.692f
C10170 VDD.n2988 VSUBS 0.0198f
C10171 VDD.n2989 VSUBS 0.814f
C10172 VDD.n2990 VSUBS 0.0198f
C10173 VDD.n2991 VSUBS 0.865f
C10174 VDD.n2992 VSUBS 0.509f
C10175 VDD.n2993 VSUBS 0.0325f
C10176 VDD.n2994 VSUBS 0.173f
C10177 VDD.n2995 VSUBS 0.183f
C10178 VDD.n2996 VSUBS 0.0112f
C10179 VDD.n2997 VSUBS 0.00362f
C10180 VDD.n2998 VSUBS 0.00794f
C10181 VDD.n2999 VSUBS 0.0033f
C10182 VDD.n3000 VSUBS 0.00126f
C10183 VDD.n3001 VSUBS 0.0355f
C10184 VDD.n3002 VSUBS 0.00496f
C10185 VDD.n3003 VSUBS 0.0059f
C10186 VDD.n3004 VSUBS 0.00189f
C10187 VDD.n3005 VSUBS 0.00153f
C10188 VDD.n3006 VSUBS 7.87e-19
C10189 VDD.n3007 VSUBS 0.00764f
C10190 VDD.n3008 VSUBS 0.00194f
C10191 VDD.t6 VSUBS 0.499f
C10192 VDD.n3009 VSUBS 0.0198f
C10193 VDD.n3010 VSUBS 0.0712f
C10194 VDD.n3011 VSUBS 0.183f
C10195 VDD.n3012 VSUBS 0.0155f
C10196 VDD.n3013 VSUBS 0.173f
C10197 VDD.n3014 VSUBS 0.509f
C10198 VDD.n3015 VSUBS 0.00639f
C10199 VDD.n3016 VSUBS 7.87e-19
C10200 VDD.n3017 VSUBS 0.00362f
C10201 VDD.n3018 VSUBS 0.00134f
C10202 VDD.n3019 VSUBS 0.00201f
C10203 VDD.n3020 VSUBS 0.00201f
C10204 VDD.n3021 VSUBS 0.00338f
C10205 VDD.n3022 VSUBS 0.0011f
C10206 VDD.n3023 VSUBS 0.00413f
C10207 VDD.n3024 VSUBS 0.00401f
C10208 VDD.n3025 VSUBS 0.00212f
C10209 VDD.n3026 VSUBS 0.00201f
C10210 VDD.n3027 VSUBS 4.72e-19
C10211 VDD.n3028 VSUBS 0.00593f
C10212 VDD.n3029 VSUBS 0.00194f
C10213 VDD.n3030 VSUBS 0.0198f
C10214 VDD.n3031 VSUBS 0.366f
C10215 VDD.n3032 VSUBS 0.183f
C10216 VDD.n3033 VSUBS 0.0155f
C10217 VDD.n3034 VSUBS 0.173f
C10218 VDD.n3035 VSUBS 0.478f
C10219 VDD.n3036 VSUBS 0.00616f
C10220 VDD.n3037 VSUBS 7.87e-19
C10221 VDD.n3038 VSUBS 0.00346f
C10222 VDD.n3039 VSUBS 0.00134f
C10223 VDD.n3040 VSUBS 0.00201f
C10224 VDD.n3041 VSUBS 0.00177f
C10225 VDD.n3042 VSUBS 0.00165f
C10226 VDD.n3043 VSUBS 0.00307f
C10227 VDD.n3044 VSUBS 0.00102f
C10228 VDD.n3045 VSUBS 8.65e-19
C10229 VDD.n3046 VSUBS 0.00458f
C10230 VDD.n3047 VSUBS 0.00537f
C10231 VDD.n3048 VSUBS 0.025f
C10232 VDD.n3049 VSUBS 0.00307f
C10233 VDD.n3050 VSUBS 0.00602f
C10234 VDD.n3051 VSUBS 0.00649f
C10235 VDD.n3052 VSUBS 0.00307f
C10236 VDD.n3053 VSUBS 0.00649f
C10237 VDD.n3054 VSUBS 0.00602f
C10238 VDD.n3055 VSUBS 0.00307f
C10239 VDD.n3056 VSUBS 0.00496f
C10240 VDD.n3057 VSUBS 0.00543f
C10241 VDD.n3058 VSUBS 0.0026f
C10242 VDD.n3059 VSUBS 0.0026f
C10243 VDD.n3060 VSUBS 0.00543f
C10244 VDD.n3061 VSUBS 0.00507f
C10245 VDD.n3062 VSUBS 0.00295f
C10246 VDD.n3063 VSUBS 0.00295f
C10247 VDD.n3064 VSUBS 0.00507f
C10248 VDD.n3065 VSUBS 0.0046f
C10249 VDD.n3066 VSUBS 0.00307f
C10250 VDD.n3067 VSUBS 0.00637f
C10251 VDD.n3068 VSUBS 0.00614f
C10252 VDD.n3069 VSUBS 0.00307f
C10253 VDD.n3070 VSUBS 0.0046f
C10254 VDD.n3071 VSUBS 0.00507f
C10255 VDD.n3072 VSUBS 0.00295f
C10256 VDD.n3073 VSUBS 0.00295f
C10257 VDD.n3074 VSUBS 0.00507f
C10258 VDD.n3075 VSUBS 0.00519f
C10259 VDD.n3076 VSUBS 0.00283f
C10260 VDD.n3077 VSUBS 0.00283f
C10261 VDD.n3078 VSUBS 0.00519f
C10262 VDD.n3079 VSUBS 0.00472f
C10263 VDD.n3080 VSUBS 0.00307f
C10264 VDD.n3081 VSUBS 0.00602f
C10265 VDD.n3082 VSUBS 0.00649f
C10266 VDD.n3083 VSUBS 0.00307f
C10267 VDD.n3084 VSUBS 0.00649f
C10268 VDD.n3085 VSUBS 0.00602f
C10269 VDD.n3086 VSUBS 0.00307f
C10270 VDD.n3087 VSUBS 0.00496f
C10271 VDD.n3088 VSUBS 0.00543f
C10272 VDD.n3089 VSUBS 0.0026f
C10273 VDD.n3090 VSUBS 0.0026f
C10274 VDD.n3091 VSUBS 0.00543f
C10275 VDD.n3092 VSUBS 0.00507f
C10276 VDD.n3093 VSUBS 0.00295f
C10277 VDD.n3094 VSUBS 0.00295f
C10278 VDD.n3095 VSUBS 0.00507f
C10279 VDD.n3096 VSUBS 0.0046f
C10280 VDD.n3097 VSUBS 0.00307f
C10281 VDD.n3098 VSUBS 0.00637f
C10282 VDD.n3099 VSUBS 0.00614f
C10283 VDD.n3100 VSUBS 0.00307f
C10284 VDD.n3101 VSUBS 0.0046f
C10285 VDD.n3102 VSUBS 0.00507f
C10286 VDD.n3103 VSUBS 0.00295f
C10287 VDD.n3104 VSUBS 0.00295f
C10288 VDD.n3105 VSUBS 0.00507f
C10289 VDD.n3106 VSUBS 0.00519f
C10290 VDD.n3107 VSUBS 0.00283f
C10291 VDD.n3108 VSUBS 0.00283f
C10292 VDD.n3109 VSUBS 0.00519f
C10293 VDD.n3110 VSUBS 0.00472f
C10294 VDD.n3111 VSUBS 0.00307f
C10295 VDD.n3112 VSUBS 0.00602f
C10296 VDD.n3113 VSUBS 0.00649f
C10297 VDD.n3114 VSUBS 0.00307f
C10298 VDD.n3115 VSUBS 0.00649f
C10299 VDD.n3116 VSUBS 0.00602f
C10300 VDD.n3117 VSUBS 0.00307f
C10301 VDD.n3118 VSUBS 0.00496f
C10302 VDD.n3119 VSUBS 0.00543f
C10303 VDD.n3120 VSUBS 0.0026f
C10304 VDD.n3121 VSUBS 0.0026f
C10305 VDD.n3122 VSUBS 0.00543f
C10306 VDD.n3123 VSUBS 0.00507f
C10307 VDD.n3124 VSUBS 0.00295f
C10308 VDD.n3125 VSUBS 0.00295f
C10309 VDD.n3126 VSUBS 0.00507f
C10310 VDD.n3127 VSUBS 0.0046f
C10311 VDD.n3128 VSUBS 0.00307f
C10312 VDD.n3129 VSUBS 0.00637f
C10313 VDD.n3130 VSUBS 0.00614f
C10314 VDD.n3131 VSUBS 0.00307f
C10315 VDD.n3132 VSUBS 0.0046f
C10316 VDD.n3133 VSUBS 0.00507f
C10317 VDD.n3134 VSUBS 0.00295f
C10318 VDD.n3135 VSUBS 0.00295f
C10319 VDD.n3136 VSUBS 0.00507f
C10320 VDD.n3137 VSUBS 0.00519f
C10321 VDD.n3138 VSUBS 0.00283f
C10322 VDD.n3139 VSUBS 0.00283f
C10323 VDD.n3140 VSUBS 0.00519f
C10324 VDD.n3141 VSUBS 0.00472f
C10325 VDD.n3142 VSUBS 0.00307f
C10326 VDD.n3143 VSUBS 0.00602f
C10327 VDD.n3144 VSUBS 0.00649f
C10328 VDD.n3145 VSUBS 0.00307f
C10329 VDD.n3146 VSUBS 0.00649f
C10330 VDD.n3147 VSUBS 0.00602f
C10331 VDD.n3148 VSUBS 0.00307f
C10332 VDD.n3149 VSUBS 0.00496f
C10333 VDD.n3150 VSUBS 0.00543f
C10334 VDD.n3151 VSUBS 0.0026f
C10335 VDD.n3152 VSUBS 0.0026f
C10336 VDD.n3153 VSUBS 0.00543f
C10337 VDD.n3154 VSUBS 0.00507f
C10338 VDD.n3155 VSUBS 0.00295f
C10339 VDD.n3156 VSUBS 0.00295f
C10340 VDD.n3157 VSUBS 0.00507f
C10341 VDD.n3158 VSUBS 0.0046f
C10342 VDD.n3159 VSUBS 0.00307f
C10343 VDD.n3160 VSUBS 0.00637f
C10344 VDD.n3161 VSUBS 0.00614f
C10345 VDD.n3162 VSUBS 0.00307f
C10346 VDD.n3163 VSUBS 0.0046f
C10347 VDD.n3164 VSUBS 0.00507f
C10348 VDD.n3165 VSUBS 0.00295f
C10349 VDD.n3166 VSUBS 0.00295f
C10350 VDD.n3167 VSUBS 0.00507f
C10351 VDD.n3168 VSUBS 0.00519f
C10352 VDD.n3169 VSUBS 0.00283f
C10353 VDD.n3170 VSUBS 0.00283f
C10354 VDD.n3171 VSUBS 0.00519f
C10355 VDD.n3172 VSUBS 0.00472f
C10356 VDD.n3173 VSUBS 0.00307f
C10357 VDD.n3174 VSUBS 0.00602f
C10358 VDD.n3175 VSUBS 0.00649f
C10359 VDD.n3176 VSUBS 0.00307f
C10360 VDD.n3177 VSUBS 0.00649f
C10361 VDD.n3178 VSUBS 0.00602f
C10362 VDD.n3179 VSUBS 0.00307f
C10363 VDD.n3180 VSUBS 0.00496f
C10364 VDD.n3181 VSUBS 0.00543f
C10365 VDD.n3182 VSUBS 0.0026f
C10366 VDD.n3183 VSUBS 0.0026f
C10367 VDD.n3184 VSUBS 0.00543f
C10368 VDD.n3185 VSUBS 0.00507f
C10369 VDD.n3186 VSUBS 0.00295f
C10370 VDD.n3187 VSUBS 0.00295f
C10371 VDD.n3188 VSUBS 0.00507f
C10372 VDD.n3189 VSUBS 0.0046f
C10373 VDD.n3190 VSUBS 0.00307f
C10374 VDD.n3191 VSUBS 0.00637f
C10375 VDD.n3192 VSUBS 0.00614f
C10376 VDD.n3193 VSUBS 0.00307f
C10377 VDD.n3194 VSUBS 0.0046f
C10378 VDD.n3195 VSUBS 0.00507f
C10379 VDD.n3196 VSUBS 0.00295f
C10380 VDD.n3197 VSUBS 0.00295f
C10381 VDD.n3198 VSUBS 0.00507f
C10382 VDD.n3199 VSUBS 0.00519f
C10383 VDD.n3200 VSUBS 0.00283f
C10384 VDD.n3201 VSUBS 0.00283f
C10385 VDD.n3202 VSUBS 0.00519f
C10386 VDD.n3203 VSUBS 0.00472f
C10387 VDD.n3204 VSUBS 0.00307f
C10388 VDD.n3205 VSUBS 0.00602f
C10389 VDD.n3206 VSUBS 0.00649f
C10390 VDD.n3207 VSUBS 0.00307f
C10391 VDD.n3208 VSUBS 0.00649f
C10392 VDD.n3209 VSUBS 0.00602f
C10393 VDD.n3210 VSUBS 0.00307f
C10394 VDD.n3211 VSUBS 0.00496f
C10395 VDD.n3212 VSUBS 0.00543f
C10396 VDD.n3213 VSUBS 0.0026f
C10397 VDD.n3214 VSUBS 0.0026f
C10398 VDD.n3215 VSUBS 0.00543f
C10399 VDD.n3216 VSUBS 0.00507f
C10400 VDD.n3217 VSUBS 0.00295f
C10401 VDD.n3218 VSUBS 0.00295f
C10402 VDD.n3219 VSUBS 0.00507f
C10403 VDD.n3220 VSUBS 0.0046f
C10404 VDD.n3221 VSUBS 0.00307f
C10405 VDD.n3222 VSUBS 0.00637f
C10406 VDD.n3223 VSUBS 0.00614f
C10407 VDD.n3224 VSUBS 0.00307f
C10408 VDD.n3225 VSUBS 0.0046f
C10409 VDD.n3226 VSUBS 0.00507f
C10410 VDD.n3227 VSUBS 0.00295f
C10411 VDD.n3228 VSUBS 0.00295f
C10412 VDD.n3229 VSUBS 0.00507f
C10413 VDD.n3230 VSUBS 0.00519f
C10414 VDD.n3231 VSUBS 0.00283f
C10415 VDD.n3232 VSUBS 0.00283f
C10416 VDD.n3233 VSUBS 0.00519f
C10417 VDD.n3234 VSUBS 0.00472f
C10418 VDD.n3235 VSUBS 0.00307f
C10419 VDD.n3236 VSUBS 0.00602f
C10420 VDD.n3237 VSUBS 0.00649f
C10421 VDD.n3238 VSUBS 0.00307f
C10422 VDD.n3239 VSUBS 0.00649f
C10423 VDD.n3240 VSUBS 0.00602f
C10424 VDD.n3241 VSUBS 0.00307f
C10425 VDD.n3242 VSUBS 0.00496f
C10426 VDD.n3243 VSUBS 0.00543f
C10427 VDD.n3244 VSUBS 0.0026f
C10428 VDD.n3245 VSUBS 0.0026f
C10429 VDD.n3246 VSUBS 0.00543f
C10430 VDD.n3247 VSUBS 0.00507f
C10431 VDD.n3248 VSUBS 0.00295f
C10432 VDD.n3249 VSUBS 0.00295f
C10433 VDD.n3250 VSUBS 0.00507f
C10434 VDD.n3251 VSUBS 0.0046f
C10435 VDD.n3252 VSUBS 0.00307f
C10436 VDD.n3253 VSUBS 0.00637f
C10437 VDD.n3254 VSUBS 0.00614f
C10438 VDD.n3255 VSUBS 0.00307f
C10439 VDD.n3256 VSUBS 0.0046f
C10440 VDD.n3257 VSUBS 0.00507f
C10441 VDD.n3258 VSUBS 0.00295f
C10442 VDD.n3259 VSUBS 0.00295f
C10443 VDD.n3260 VSUBS 0.00507f
C10444 VDD.n3261 VSUBS 0.00519f
C10445 VDD.n3262 VSUBS 0.00283f
C10446 VDD.n3263 VSUBS 0.00283f
C10447 VDD.n3264 VSUBS 0.00519f
C10448 VDD.n3265 VSUBS 0.00472f
C10449 VDD.n3266 VSUBS 0.00307f
C10450 VDD.n3267 VSUBS 0.00602f
C10451 VDD.n3268 VSUBS 0.00649f
C10452 VDD.n3269 VSUBS 0.00307f
C10453 VDD.n3270 VSUBS 0.00649f
C10454 VDD.n3271 VSUBS 0.00602f
C10455 VDD.n3272 VSUBS 0.00307f
C10456 VDD.n3273 VSUBS 0.00496f
C10457 VDD.n3274 VSUBS 0.00543f
C10458 VDD.n3275 VSUBS 0.0026f
C10459 VDD.n3276 VSUBS 0.0026f
C10460 VDD.n3277 VSUBS 0.00543f
C10461 VDD.n3278 VSUBS 0.00507f
C10462 VDD.n3279 VSUBS 0.00295f
C10463 VDD.n3280 VSUBS 0.00295f
C10464 VDD.n3281 VSUBS 0.00507f
C10465 VDD.n3282 VSUBS 0.0046f
C10466 VDD.n3283 VSUBS 0.00307f
C10467 VDD.n3284 VSUBS 0.00637f
C10468 VDD.n3285 VSUBS 0.00614f
C10469 VDD.n3286 VSUBS 0.00307f
C10470 VDD.n3287 VSUBS 0.0046f
C10471 VDD.n3288 VSUBS 0.00507f
C10472 VDD.n3289 VSUBS 0.00295f
C10473 VDD.n3290 VSUBS 0.00295f
C10474 VDD.n3291 VSUBS 0.00507f
C10475 VDD.n3292 VSUBS 0.00519f
C10476 VDD.n3293 VSUBS 0.00283f
C10477 VDD.n3294 VSUBS 0.00283f
C10478 VDD.n3295 VSUBS 0.00519f
C10479 VDD.n3296 VSUBS 0.00472f
C10480 VDD.n3297 VSUBS 0.00307f
C10481 VDD.n3298 VSUBS 0.00602f
C10482 VDD.n3299 VSUBS 0.00649f
C10483 VDD.n3300 VSUBS 0.00307f
C10484 VDD.n3301 VSUBS 0.00649f
C10485 VDD.n3302 VSUBS 0.00602f
C10486 VDD.n3303 VSUBS 0.00307f
C10487 VDD.n3304 VSUBS 0.00496f
C10488 VDD.n3305 VSUBS 0.00543f
C10489 VDD.n3306 VSUBS 0.0026f
C10490 VDD.n3307 VSUBS 0.0026f
C10491 VDD.n3308 VSUBS 0.00543f
C10492 VDD.n3309 VSUBS 0.00507f
C10493 VDD.n3310 VSUBS 0.00295f
C10494 VDD.n3311 VSUBS 0.00295f
C10495 VDD.n3312 VSUBS 0.00507f
C10496 VDD.n3313 VSUBS 0.0046f
C10497 VDD.n3314 VSUBS 0.00307f
C10498 VDD.n3315 VSUBS 0.00637f
C10499 VDD.n3316 VSUBS 0.00614f
C10500 VDD.n3317 VSUBS 0.00307f
C10501 VDD.n3318 VSUBS 0.0046f
C10502 VDD.n3319 VSUBS 0.00507f
C10503 VDD.n3320 VSUBS 0.00295f
C10504 VDD.n3321 VSUBS 0.00295f
C10505 VDD.n3322 VSUBS 0.00507f
C10506 VDD.n3323 VSUBS 0.00519f
C10507 VDD.n3324 VSUBS 0.00283f
C10508 VDD.n3325 VSUBS 0.00283f
C10509 VDD.n3326 VSUBS 0.00519f
C10510 VDD.n3327 VSUBS 0.00472f
C10511 VDD.n3328 VSUBS 0.00307f
C10512 VDD.n3329 VSUBS 0.00602f
C10513 VDD.n3330 VSUBS 0.00649f
C10514 VDD.n3331 VSUBS 0.00307f
C10515 VDD.n3332 VSUBS 0.00649f
C10516 VDD.n3333 VSUBS 0.00602f
C10517 VDD.n3334 VSUBS 0.00307f
C10518 VDD.n3335 VSUBS 0.00496f
C10519 VDD.n3336 VSUBS 0.00543f
C10520 VDD.n3337 VSUBS 0.0026f
C10521 VDD.n3338 VSUBS 0.0026f
C10522 VDD.n3339 VSUBS 0.00543f
C10523 VDD.n3340 VSUBS 0.00507f
C10524 VDD.n3341 VSUBS 0.00295f
C10525 VDD.n3342 VSUBS 0.00295f
C10526 VDD.n3343 VSUBS 0.00507f
C10527 VDD.n3344 VSUBS 0.0046f
C10528 VDD.n3345 VSUBS 0.00307f
C10529 VDD.n3346 VSUBS 0.00637f
C10530 VDD.n3347 VSUBS 0.00614f
C10531 VDD.n3348 VSUBS 0.00307f
C10532 VDD.n3349 VSUBS 0.0046f
C10533 VDD.n3350 VSUBS 0.00507f
C10534 VDD.n3351 VSUBS 0.00295f
C10535 VDD.n3352 VSUBS 0.00295f
C10536 VDD.n3353 VSUBS 0.00507f
C10537 VDD.n3354 VSUBS 0.00519f
C10538 VDD.n3355 VSUBS 0.00283f
C10539 VDD.n3356 VSUBS 0.00283f
C10540 VDD.n3357 VSUBS 0.00519f
C10541 VDD.n3358 VSUBS 0.00472f
C10542 VDD.n3359 VSUBS 0.00307f
C10543 VDD.n3360 VSUBS 0.00602f
C10544 VDD.n3361 VSUBS 0.00649f
C10545 VDD.n3362 VSUBS 0.00307f
C10546 VDD.n3363 VSUBS 0.00649f
C10547 VDD.n3364 VSUBS 0.00602f
C10548 VDD.n3365 VSUBS 0.00307f
C10549 VDD.n3366 VSUBS 0.00496f
C10550 VDD.n3367 VSUBS 0.00543f
C10551 VDD.n3368 VSUBS 0.0026f
C10552 VDD.n3369 VSUBS 0.0026f
C10553 VDD.n3370 VSUBS 0.00543f
C10554 VDD.n3371 VSUBS 0.00507f
C10555 VDD.n3372 VSUBS 0.00295f
C10556 VDD.n3373 VSUBS 0.00295f
C10557 VDD.n3374 VSUBS 0.00507f
C10558 VDD.n3375 VSUBS 0.0046f
C10559 VDD.n3376 VSUBS 0.00307f
C10560 VDD.n3377 VSUBS 0.00637f
C10561 VDD.n3378 VSUBS 0.00614f
C10562 VDD.n3379 VSUBS 0.00307f
C10563 VDD.n3380 VSUBS 0.0046f
C10564 VDD.n3381 VSUBS 0.00507f
C10565 VDD.n3382 VSUBS 0.00295f
C10566 VDD.n3383 VSUBS 0.00295f
C10567 VDD.n3384 VSUBS 0.00507f
C10568 VDD.n3385 VSUBS 0.00519f
C10569 VDD.n3386 VSUBS 0.00283f
C10570 VDD.n3387 VSUBS 0.00283f
C10571 VDD.n3388 VSUBS 0.00519f
C10572 VDD.n3389 VSUBS 0.00472f
C10573 VDD.n3390 VSUBS 0.00378f
C10574 VDD.n3391 VSUBS 0.00134f
C10575 VDD.n3392 VSUBS 0.00741f
C10576 VDD.n3393 VSUBS 0.00194f
C10577 VDD.n3394 VSUBS 0.0198f
C10578 VDD.n3395 VSUBS 0.539f
C10579 VDD.n3396 VSUBS 0.183f
C10580 VDD.n3397 VSUBS 0.0155f
C10581 VDD.n3398 VSUBS 0.173f
C10582 VDD.n3399 VSUBS 0.509f
C10583 VDD.n3400 VSUBS 0.00661f
C10584 VDD.n3401 VSUBS 7.87e-19
C10585 VDD.n3402 VSUBS 0.00378f
C10586 VDD.n3403 VSUBS 0.00134f
C10587 VDD.n3404 VSUBS 0.00165f
C10588 VDD.n3405 VSUBS 0.00142f
C10589 VDD.n3406 VSUBS 0.00201f
C10590 VDD.n3407 VSUBS 0.0046f
C10591 VDD.n3408 VSUBS 0.0046f
C10592 VDD.n3409 VSUBS 0.00248f
C10593 VDD.n3410 VSUBS 0.00362f
C10594 VDD.n3411 VSUBS 0.00134f
C10595 VDD.n3412 VSUBS 0.00719f
C10596 VDD.n3413 VSUBS 0.00194f
C10597 VDD.n3414 VSUBS 0.0198f
C10598 VDD.n3415 VSUBS 0.539f
C10599 VDD.n3416 VSUBS 0.183f
C10600 VDD.n3417 VSUBS 0.0155f
C10601 VDD.n3418 VSUBS 0.112f
C10602 VDD.t61 VSUBS 0.0712f
C10603 VDD.n3419 VSUBS 0.499f
C10604 VDD.n3420 VSUBS 0.00684f
C10605 VDD.n3421 VSUBS 0.0011f
C10606 VDD.n3422 VSUBS 0.00362f
C10607 VDD.n3423 VSUBS 0.00134f
C10608 VDD.n3424 VSUBS 9.44e-19
C10609 VDD.n3425 VSUBS 0.00118f
C10610 VDD.n3426 VSUBS 0.00248f
C10611 VDD.n3427 VSUBS 0.00437f
C10612 VDD.n3428 VSUBS 0.00484f
C10613 VDD.n3429 VSUBS 0.00212f
C10614 VDD.n3430 VSUBS 0.00106f
C10615 VDD.n3431 VSUBS 0.00346f
C10616 VDD.n3432 VSUBS 0.00134f
C10617 VDD.n3433 VSUBS 0.00696f
C10618 VDD.n3434 VSUBS 0.00194f
C10619 VDD.n3435 VSUBS 0.0198f
C10620 VDD.n3436 VSUBS 0.539f
C10621 VDD.n3437 VSUBS 0.183f
C10622 VDD.n3438 VSUBS 0.0155f
C10623 VDD.n3439 VSUBS 0.173f
C10624 VDD.n3440 VSUBS 0.509f
C10625 VDD.n3441 VSUBS 0.00707f
C10626 VDD.n3442 VSUBS 0.00142f
C10627 VDD.n3443 VSUBS 0.00346f
C10628 VDD.n3444 VSUBS 0.00134f
C10629 VDD.n3445 VSUBS 0.00177f
C10630 VDD.n3446 VSUBS 0.00212f
C10631 VDD.n3447 VSUBS 0.00413f
C10632 VDD.n3448 VSUBS 0.0046f
C10633 VDD.n3449 VSUBS 0.00212f
C10634 VDD.n3450 VSUBS 0.00142f
C10635 VDD.n3451 VSUBS 0.0033f
C10636 VDD.n3452 VSUBS 0.00134f
C10637 VDD.n3453 VSUBS 0.00673f
C10638 VDD.n3454 VSUBS 0.00194f
C10639 VDD.n3455 VSUBS 0.0198f
C10640 VDD.n3456 VSUBS 0.539f
C10641 VDD.n3457 VSUBS 0.183f
C10642 VDD.n3458 VSUBS 0.0155f
C10643 VDD.n3459 VSUBS 0.173f
C10644 VDD.t42 VSUBS 0.397f
C10645 VDD.n3460 VSUBS 0.234f
C10646 VDD.n3461 VSUBS 0.0073f
C10647 VDD.n3462 VSUBS 0.00149f
C10648 VDD.n3463 VSUBS 0.00134f
C10649 VDD.n3464 VSUBS 0.00134f
C10650 VDD.n3465 VSUBS 0.00201f
C10651 VDD.n3466 VSUBS 0.00201f
C10652 VDD.n3467 VSUBS 0.00283f
C10653 VDD.n3468 VSUBS 0.00389f
C10654 VDD.n3469 VSUBS 0.00413f
C10655 VDD.n3470 VSUBS 0.00236f
C10656 VDD.n3471 VSUBS 0.00189f
C10657 VDD.n3472 VSUBS 0.00252f
C10658 VDD.n3473 VSUBS 0.00134f
C10659 VDD.n3474 VSUBS 0.0065f
C10660 VDD.n3475 VSUBS 0.00194f
C10661 VDD.n3476 VSUBS 0.0198f
C10662 VDD.n3477 VSUBS 0.417f
C10663 VDD.n3478 VSUBS 0.183f
C10664 VDD.n3479 VSUBS 0.0155f
C10665 VDD.n3480 VSUBS 0.173f
C10666 VDD.n3481 VSUBS 0.509f
C10667 VDD.n3482 VSUBS 0.00753f
C10668 VDD.n3483 VSUBS 0.00149f
C10669 VDD.n3484 VSUBS 0.00126f
C10670 VDD.n3485 VSUBS 0.00134f
C10671 VDD.n3486 VSUBS 0.00201f
C10672 VDD.n3487 VSUBS 0.00189f
C10673 VDD.n3488 VSUBS 0.00142f
C10674 VDD.n3489 VSUBS 9.44e-19
C10675 VDD.n3490 VSUBS 0.00244f
C10676 VDD.n3491 VSUBS 0.00319f
C10677 VDD.n3492 VSUBS 0.00295f
C10678 VDD.n3493 VSUBS 0.00248f
C10679 VDD.n3494 VSUBS 0.00236f
C10680 VDD.n3495 VSUBS 0.00205f
C10681 VDD.n3496 VSUBS 0.00134f
C10682 VDD.n3497 VSUBS 0.00627f
C10683 VDD.n3498 VSUBS 0.00194f
C10684 VDD.n3499 VSUBS 0.0198f
C10685 VDD.n3500 VSUBS 0.539f
C10686 VDD.n3501 VSUBS 0.183f
C10687 VDD.n3502 VSUBS 0.0155f
C10688 VDD.n3503 VSUBS 0.173f
C10689 VDD.n3504 VSUBS 0.0155f
C10690 VDD.n3505 VSUBS 0.692f
C10691 VDD.n3506 VSUBS 0.0198f
C10692 VDD.n3507 VSUBS 0.234f
C10693 VDD.t45 VSUBS 0.356f
C10694 VDD.n3508 VSUBS 0.458f
C10695 VDD.n3509 VSUBS 0.00776f
C10696 VDD.n3510 VSUBS 0.00149f
C10697 VDD.n3511 VSUBS 0.00126f
C10698 VDD.n3512 VSUBS 0.00189f
C10699 VDD.n3513 VSUBS 0.00153f
C10700 VDD.n3514 VSUBS 0.0013f
C10701 VDD.n3515 VSUBS 0.00102f
C10702 VDD.n3516 VSUBS 8.65e-19
C10703 VDD.n3517 VSUBS 0.00283f
C10704 VDD.n3518 VSUBS 0.00366f
C10705 VDD.n3519 VSUBS 0.00283f
C10706 VDD.n3520 VSUBS 0.00283f
C10707 VDD.n3521 VSUBS 0.0138f
C10708 VDD.n3522 VSUBS 0.00354f
C10709 VDD.n3523 VSUBS 0.00118f
C10710 VDD.n3524 VSUBS 0.00212f
C10711 VDD.n3525 VSUBS 0.00342f
C10712 VDD.n3526 VSUBS 0.00177f
C10713 VDD.n3527 VSUBS 0.00177f
C10714 VDD.n3528 VSUBS 0.00118f
C10715 VDD.n3529 VSUBS 0.0138f
C10716 VDD.n3530 VSUBS 0.00401f
C10717 VDD.n3531 VSUBS 0.00267f
C10718 VDD.n3532 VSUBS 0.00295f
C10719 VDD.n3533 VSUBS 0.00307f
C10720 VDD.n3534 VSUBS 0.00401f
C10721 VDD.n3535 VSUBS 0.00283f
C10722 VDD.n3536 VSUBS 0.00425f
C10723 VDD.n3537 VSUBS 0.00201f
C10724 VDD.n3538 VSUBS 0.00134f
C10725 VDD.n3539 VSUBS 0.00299f
C10726 VDD.n3540 VSUBS 0.00134f
C10727 VDD.n3541 VSUBS 0.00627f
C10728 VDD.n3542 VSUBS 0.00194f
C10729 VDD.n3543 VSUBS 0.0198f
C10730 VDD.n3544 VSUBS 0.692f
C10731 VDD.n3545 VSUBS 0.0155f
C10732 VDD.n3546 VSUBS 0.692f
C10733 VDD.n3547 VSUBS 0.0198f
C10734 VDD.n3548 VSUBS 0.539f
C10735 VDD.n3549 VSUBS 0.509f
C10736 VDD.n3550 VSUBS 0.0155f
C10737 VDD.n3551 VSUBS 0.0305f
C10738 VDD.t88 VSUBS 0.153f
C10739 VDD.n3552 VSUBS 0.173f
C10740 VDD.n3553 VSUBS 0.00776f
C10741 VDD.n3554 VSUBS 0.00205f
C10742 VDD.n3555 VSUBS 0.00134f
C10743 VDD.n3556 VSUBS 0.00201f
C10744 VDD.n3557 VSUBS 0.00153f
C10745 VDD.n3558 VSUBS 0.00177f
C10746 VDD.n3559 VSUBS 0.00602f
C10747 VDD.n3560 VSUBS 0.00496f
C10748 VDD.n3561 VSUBS 0.00315f
C10749 VDD.n3562 VSUBS 0.00315f
C10750 VDD.n3563 VSUBS 0.00134f
C10751 VDD.n3564 VSUBS 0.0065f
C10752 VDD.n3565 VSUBS 0.00194f
C10753 VDD.n3566 VSUBS 0.0198f
C10754 VDD.n3567 VSUBS 0.539f
C10755 VDD.n3568 VSUBS 0.509f
C10756 VDD.n3569 VSUBS 0.0155f
C10757 VDD.n3570 VSUBS 0.173f
C10758 VDD.n3571 VSUBS 0.183f
C10759 VDD.n3572 VSUBS 0.00753f
C10760 VDD.n3573 VSUBS 0.00205f
C10761 VDD.n3574 VSUBS 0.00134f
C10762 VDD.n3575 VSUBS 0.00153f
C10763 VDD.n3576 VSUBS 0.00153f
C10764 VDD.n3577 VSUBS 0.00201f
C10765 VDD.n3578 VSUBS 0.00448f
C10766 VDD.n3579 VSUBS 0.00472f
C10767 VDD.n3580 VSUBS 0.00248f
C10768 VDD.n3581 VSUBS 0.0033f
C10769 VDD.n3582 VSUBS 0.0033f
C10770 VDD.n3583 VSUBS 0.00134f
C10771 VDD.n3584 VSUBS 0.00673f
C10772 VDD.n3585 VSUBS 0.00194f
C10773 VDD.n3586 VSUBS 0.0198f
C10774 VDD.n3587 VSUBS 0.539f
C10775 VDD.t29 VSUBS 0.448f
C10776 VDD.n3588 VSUBS 0.214f
C10777 VDD.n3589 VSUBS 0.0155f
C10778 VDD.n3590 VSUBS 0.173f
C10779 VDD.n3591 VSUBS 0.183f
C10780 VDD.n3592 VSUBS 0.0073f
C10781 VDD.n3593 VSUBS 0.00173f
C10782 VDD.n3594 VSUBS 0.00134f
C10783 VDD.n3595 VSUBS 8.26e-19
C10784 VDD.n3596 VSUBS 0.0013f
C10785 VDD.n3597 VSUBS 0.00248f
C10786 VDD.n3598 VSUBS 0.00425f
C10787 VDD.n3599 VSUBS 0.00496f
C10788 VDD.n3600 VSUBS 0.00212f
C10789 VDD.n3601 VSUBS 9.44e-19
C10790 VDD.n3602 VSUBS 0.00346f
C10791 VDD.n3603 VSUBS 0.00346f
C10792 VDD.n3604 VSUBS 0.00134f
C10793 VDD.n3605 VSUBS 0.00696f
C10794 VDD.n3606 VSUBS 0.00194f
C10795 VDD.n3607 VSUBS 0.0198f
C10796 VDD.n3608 VSUBS 0.387f
C10797 VDD.n3609 VSUBS 0.509f
C10798 VDD.n3610 VSUBS 0.0155f
C10799 VDD.n3611 VSUBS 0.173f
C10800 VDD.n3612 VSUBS 0.183f
C10801 VDD.n3613 VSUBS 0.00707f
C10802 VDD.n3614 VSUBS 0.00142f
C10803 VDD.n3615 VSUBS 0.00134f
C10804 VDD.n3616 VSUBS 0.00189f
C10805 VDD.n3617 VSUBS 0.00212f
C10806 VDD.n3618 VSUBS 0.00401f
C10807 VDD.n3619 VSUBS 0.0046f
C10808 VDD.n3620 VSUBS 0.00224f
C10809 VDD.n3621 VSUBS 0.00142f
C10810 VDD.n3622 VSUBS 0.00338f
C10811 VDD.n3623 VSUBS 0.00719f
C10812 VDD.n3624 VSUBS 0.00194f
C10813 VDD.n3625 VSUBS 0.0198f
C10814 VDD.n3626 VSUBS 0.539f
C10815 VDD.n3627 VSUBS 0.438f
C10816 VDD.n3628 VSUBS 0.0155f
C10817 VDD.n3629 VSUBS 0.173f
C10818 VDD.n3630 VSUBS 0.183f
C10819 VDD.n3631 VSUBS 0.00684f
C10820 VDD.n3632 VSUBS 0.00134f
C10821 VDD.n3633 VSUBS 0.00134f
C10822 VDD.n3634 VSUBS 0.00201f
C10823 VDD.n3635 VSUBS 0.00201f
C10824 VDD.n3636 VSUBS 0.00362f
C10825 VDD.n3637 VSUBS 0.00134f
C10826 VDD.n3638 VSUBS 0.00378f
C10827 VDD.n3639 VSUBS 0.00413f
C10828 VDD.n3640 VSUBS 0.00248f
C10829 VDD.n3641 VSUBS 0.00189f
C10830 VDD.n3642 VSUBS 0.00322f
C10831 VDD.n3643 VSUBS 0.00134f
C10832 VDD.n3644 VSUBS 0.00201f
C10833 VDD.n3645 VSUBS 0.00189f
C10834 VDD.n3646 VSUBS 0.0013f
C10835 VDD.n3647 VSUBS 0.00741f
C10836 VDD.n3648 VSUBS 0.00194f
C10837 VDD.t17 VSUBS 0.407f
C10838 VDD.n3649 VSUBS 0.0198f
C10839 VDD.n3650 VSUBS 0.204f
C10840 VDD.n3651 VSUBS 0.509f
C10841 VDD.n3652 VSUBS 0.0155f
C10842 VDD.n3653 VSUBS 0.173f
C10843 VDD.n3654 VSUBS 0.183f
C10844 VDD.n3655 VSUBS 0.00661f
C10845 VDD.n3656 VSUBS 0.00126f
C10846 VDD.n3657 VSUBS 3.93e-19
C10847 VDD.n3658 VSUBS 5.51e-19
C10848 VDD.n3659 VSUBS 0.0033f
C10849 VDD.n3660 VSUBS 9.44e-19
C10850 VDD.n3661 VSUBS 0.00319f
C10851 VDD.n3662 VSUBS 0.00295f
C10852 VDD.n3663 VSUBS 0.0026f
C10853 VDD.n3664 VSUBS 0.00236f
C10854 VDD.n3665 VSUBS 0.00307f
C10855 VDD.n3666 VSUBS 0.00118f
C10856 VDD.n3667 VSUBS 0.00177f
C10857 VDD.n3668 VSUBS 0.00165f
C10858 VDD.n3669 VSUBS 0.0013f
C10859 VDD.n3670 VSUBS 0.0011f
C10860 VDD.n3671 VSUBS 0.00764f
C10861 VDD.n3672 VSUBS 0.00194f
C10862 VDD.n3673 VSUBS 0.0198f
C10863 VDD.n3674 VSUBS 0.539f
C10864 VDD.n3675 VSUBS 0.509f
C10865 VDD.n3676 VSUBS 0.0155f
C10866 VDD.n3677 VSUBS 0.173f
C10867 VDD.n3678 VSUBS 0.183f
C10868 VDD.n3679 VSUBS 0.00639f
C10869 VDD.n3680 VSUBS 3.93e-19
C10870 VDD.n3681 VSUBS 7.08e-19
C10871 VDD.n3682 VSUBS 0.00346f
C10872 VDD.n3683 VSUBS 0.0011f
C10873 VDD.n3684 VSUBS 0.00354f
C10874 VDD.n3685 VSUBS 0.00283f
C10875 VDD.n3686 VSUBS 0.00271f
C10876 VDD.n3687 VSUBS 0.00248f
C10877 VDD.n3688 VSUBS 0.00291f
C10878 VDD.n3689 VSUBS 0.00126f
C10879 VDD.n3690 VSUBS 7.08e-19
C10880 VDD.n3691 VSUBS 0.00106f
C10881 VDD.n3692 VSUBS 0.00189f
C10882 VDD.n3693 VSUBS 0.00177f
C10883 VDD.n3694 VSUBS 0.00593f
C10884 VDD.n3695 VSUBS 0.00194f
C10885 VDD.n3696 VSUBS 0.0198f
C10886 VDD.n3697 VSUBS 0.519f
C10887 VDD.t143 VSUBS 0.173f
C10888 VDD.n3698 VSUBS 0.509f
C10889 VDD.n3699 VSUBS 0.0155f
C10890 VDD.n3700 VSUBS 0.173f
C10891 VDD.n3701 VSUBS 0.0305f
C10892 VDD.n3702 VSUBS 0.00616f
C10893 VDD.n3703 VSUBS 7.08e-19
C10894 VDD.n3704 VSUBS 5.51e-19
C10895 VDD.n3705 VSUBS 0.00362f
C10896 VDD.n3706 VSUBS 0.00126f
C10897 VDD.n3707 VSUBS 0.00283f
C10898 VDD.n3708 VSUBS 0.00307f
C10899 VDD.n3709 VSUBS 0.00401f
C10900 VDD.n3710 VSUBS 0.00322f
C10901 VDD.n3711 VSUBS 0.00126f
C10902 VDD.n3712 VSUBS 0.00437f
C10903 VDD.n3713 VSUBS 0.00201f
C10904 VDD.n3714 VSUBS 9.44e-19
C10905 VDD.n3715 VSUBS 0.00593f
C10906 VDD.n3716 VSUBS 0.00194f
C10907 VDD.n3717 VSUBS 0.0198f
C10908 VDD.n3718 VSUBS 0.366f
C10909 VDD.n3719 VSUBS 0.183f
C10910 VDD.n3720 VSUBS 0.0155f
C10911 VDD.n3721 VSUBS 0.173f
C10912 VDD.n3722 VSUBS 0.509f
C10913 VDD.n3723 VSUBS 0.00616f
C10914 VDD.n3724 VSUBS 4.72e-19
C10915 VDD.n3725 VSUBS 0.00378f
C10916 VDD.n3726 VSUBS 0.00134f
C10917 VDD.n3727 VSUBS 0.00201f
C10918 VDD.n3728 VSUBS 0.00153f
C10919 VDD.n3729 VSUBS 0.00165f
C10920 VDD.n3730 VSUBS 0.00614f
C10921 VDD.n3731 VSUBS 0.00496f
C10922 VDD.n3732 VSUBS 0.00393f
C10923 VDD.n3733 VSUBS 0.00134f
C10924 VDD.n3734 VSUBS 0.00764f
C10925 VDD.n3735 VSUBS 0.00194f
C10926 VDD.n3736 VSUBS 0.0198f
C10927 VDD.n3737 VSUBS 0.539f
C10928 VDD.n3738 VSUBS 0.183f
C10929 VDD.n3739 VSUBS 0.0155f
C10930 VDD.n3740 VSUBS 0.173f
C10931 VDD.t80 VSUBS 0.478f
C10932 VDD.n3741 VSUBS 0.193f
C10933 VDD.n3742 VSUBS 0.00639f
C10934 VDD.n3743 VSUBS 4.72e-19
C10935 VDD.n3744 VSUBS 0.00393f
C10936 VDD.n3745 VSUBS 0.00134f
C10937 VDD.n3746 VSUBS 0.00142f
C10938 VDD.n3747 VSUBS 0.00165f
C10939 VDD.n3748 VSUBS 0.00201f
C10940 VDD.n3749 VSUBS 0.00437f
C10941 VDD.n3750 VSUBS 0.00484f
C10942 VDD.n3751 VSUBS 0.00248f
C10943 VDD.n3752 VSUBS 0.00378f
C10944 VDD.n3753 VSUBS 0.00134f
C10945 VDD.n3754 VSUBS 0.00741f
C10946 VDD.n3755 VSUBS 0.00194f
C10947 VDD.n3756 VSUBS 0.0198f
C10948 VDD.n3757 VSUBS 0.377f
C10949 VDD.n3758 VSUBS 0.183f
C10950 VDD.n3759 VSUBS 0.0155f
C10951 VDD.n3760 VSUBS 0.173f
C10952 VDD.n3761 VSUBS 0.509f
C10953 VDD.n3762 VSUBS 0.00661f
C10954 VDD.n3763 VSUBS 7.87e-19
C10955 VDD.n3764 VSUBS 0.00378f
C10956 VDD.n3765 VSUBS 0.00134f
C10957 VDD.n3766 VSUBS 7.08e-19
C10958 VDD.n3767 VSUBS 0.00142f
C10959 VDD.n3768 VSUBS 0.00248f
C10960 VDD.n3769 VSUBS 0.00413f
C10961 VDD.n3770 VSUBS 0.00507f
C10962 VDD.n3771 VSUBS 0.00295f
C10963 VDD.n3772 VSUBS 0.00362f
C10964 VDD.n3773 VSUBS 0.00134f
C10965 VDD.n3774 VSUBS 0.00719f
C10966 VDD.n3775 VSUBS 0.00194f
C10967 VDD.n3776 VSUBS 0.0198f
C10968 VDD.n3777 VSUBS 0.539f
C10969 VDD.n3778 VSUBS 0.183f
C10970 VDD.n3779 VSUBS 0.0155f
C10971 VDD.n3780 VSUBS 0.173f
C10972 VDD.n3781 VSUBS 0.417f
C10973 VDD.n3782 VSUBS 0.00684f
C10974 VDD.n3783 VSUBS 0.0011f
C10975 VDD.n3784 VSUBS 0.00362f
C10976 VDD.n3785 VSUBS 0.00134f
C10977 VDD.n3786 VSUBS 0.00201f
C10978 VDD.n3787 VSUBS 0.00212f
C10979 VDD.n3788 VSUBS 0.00389f
C10980 VDD.n3789 VSUBS 0.0046f
C10981 VDD.n3790 VSUBS 0.00236f
C10982 VDD.n3791 VSUBS 0.00142f
C10983 VDD.n3792 VSUBS 0.00346f
C10984 VDD.n3793 VSUBS 0.00134f
C10985 VDD.n3794 VSUBS 0.00696f
C10986 VDD.n3795 VSUBS 0.00194f
C10987 VDD.t4 VSUBS 0.438f
C10988 VDD.n3796 VSUBS 0.0198f
C10989 VDD.n3797 VSUBS 0.193f
C10990 VDD.n3798 VSUBS 0.183f
C10991 VDD.n3799 VSUBS 0.0155f
C10992 VDD.n3800 VSUBS 0.173f
C10993 VDD.n3801 VSUBS 0.509f
C10994 VDD.n3802 VSUBS 0.00707f
C10995 VDD.n3803 VSUBS 0.00118f
C10996 VDD.n3804 VSUBS 0.00134f
C10997 VDD.n3805 VSUBS 0.00134f
C10998 VDD.n3806 VSUBS 0.00201f
C10999 VDD.n3807 VSUBS 0.00201f
C11000 VDD.n3808 VSUBS 0.00283f
C11001 VDD.n3809 VSUBS 0.00366f
C11002 VDD.n3810 VSUBS 0.00413f
C11003 VDD.n3811 VSUBS 0.0026f
C11004 VDD.n3812 VSUBS 0.00189f
C11005 VDD.n3813 VSUBS 0.00283f
C11006 VDD.n3814 VSUBS 0.00134f
C11007 VDD.n3815 VSUBS 0.00673f
C11008 VDD.n3816 VSUBS 0.00194f
C11009 VDD.n3817 VSUBS 0.0198f
C11010 VDD.n3818 VSUBS 0.539f
C11011 VDD.n3819 VSUBS 0.183f
C11012 VDD.n3820 VSUBS 0.0155f
C11013 VDD.n3821 VSUBS 0.173f
C11014 VDD.n3822 VSUBS 0.509f
C11015 VDD.n3823 VSUBS 0.0073f
C11016 VDD.n3824 VSUBS 0.00118f
C11017 VDD.n3825 VSUBS 0.00134f
C11018 VDD.n3826 VSUBS 0.00201f
C11019 VDD.n3827 VSUBS 0.00189f
C11020 VDD.n3828 VSUBS 0.00118f
C11021 VDD.n3829 VSUBS 0.00126f
C11022 VDD.n3830 VSUBS 7.87e-19
C11023 VDD.n3831 VSUBS 0.0026f
C11024 VDD.n3832 VSUBS 0.00319f
C11025 VDD.n3833 VSUBS 0.00295f
C11026 VDD.n3834 VSUBS 0.00271f
C11027 VDD.n3835 VSUBS 0.00236f
C11028 VDD.n3836 VSUBS 0.00236f
C11029 VDD.n3837 VSUBS 0.00134f
C11030 VDD.n3838 VSUBS 0.0065f
C11031 VDD.n3839 VSUBS 0.00194f
C11032 VDD.n3840 VSUBS 0.0198f
C11033 VDD.n3841 VSUBS 0.529f
C11034 VDD.t0 VSUBS 0.142f
C11035 VDD.n3842 VSUBS 0.0509f
C11036 VDD.n3843 VSUBS 0.0155f
C11037 VDD.n3844 VSUBS 0.173f
C11038 VDD.n3845 VSUBS 0.509f
C11039 VDD.n3846 VSUBS 0.00753f
C11040 VDD.n3847 VSUBS 0.00118f
C11041 VDD.n3848 VSUBS 0.0011f
C11042 VDD.n3849 VSUBS 0.00165f
C11043 VDD.n3850 VSUBS 0.00177f
C11044 VDD.n3851 VSUBS 0.0013f
C11045 VDD.n3852 VSUBS 0.00118f
C11046 VDD.n3853 VSUBS 8.65e-19
C11047 VDD.n3854 VSUBS 0.00283f
C11048 VDD.n3855 VSUBS 0.00342f
C11049 VDD.n3856 VSUBS 0.00283f
C11050 VDD.n3857 VSUBS 0.00283f
C11051 VDD.n3858 VSUBS 0.00236f
C11052 VDD.n3859 VSUBS 0.00134f
C11053 VDD.n3860 VSUBS 0.00134f
C11054 VDD.n3861 VSUBS 0.00627f
C11055 VDD.n3862 VSUBS 0.00194f
C11056 VDD.n3863 VSUBS 0.0198f
C11057 VDD.n3864 VSUBS 0.539f
C11058 VDD.n3865 VSUBS 0.183f
C11059 VDD.n3866 VSUBS 0.0155f
C11060 VDD.n3867 VSUBS 0.173f
C11061 VDD.n3868 VSUBS 0.0198f
C11062 VDD.n3869 VSUBS 0.519f
C11063 VDD.t19 VSUBS 0.509f
C11064 VDD.n3870 VSUBS 0.0155f
C11065 VDD.n3871 VSUBS 0.356f
C11066 VDD.n3872 VSUBS 0.0198f
C11067 VDD.n3873 VSUBS 0.539f
C11068 VDD.n3874 VSUBS 0.509f
C11069 VDD.n3875 VSUBS 0.00776f
C11070 VDD.n3876 VSUBS 0.00181f
C11071 VDD.n3877 VSUBS 0.00342f
C11072 VDD.n3878 VSUBS 0.00201f
C11073 VDD.n3879 VSUBS 0.00177f
C11074 VDD.n3880 VSUBS 0.00118f
C11075 VDD.n3881 VSUBS 0.0138f
C11076 VDD.n3882 VSUBS 0.00401f
C11077 VDD.n3883 VSUBS 0.00283f
C11078 VDD.n3884 VSUBS 0.00271f
C11079 VDD.n3885 VSUBS 0.00307f
C11080 VDD.n3886 VSUBS 0.00401f
C11081 VDD.n3887 VSUBS 0.00267f
C11082 VDD.n3888 VSUBS 0.00448f
C11083 VDD.n3889 VSUBS 0.00201f
C11084 VDD.n3890 VSUBS 0.00134f
C11085 VDD.n3891 VSUBS 0.0138f
C11086 VDD.n3892 VSUBS 0.00519f
C11087 VDD.n3893 VSUBS 0.00267f
C11088 VDD.n3894 VSUBS 0.00201f
C11089 VDD.n3895 VSUBS 0.00307f
C11090 VDD.n3896 VSUBS 0.00625f
C11091 VDD.n3897 VSUBS 0.00496f
C11092 VDD.n3898 VSUBS 0.00299f
C11093 VDD.n3899 VSUBS 0.00134f
C11094 VDD.n3900 VSUBS 0.0013f
C11095 VDD.n3901 VSUBS 0.00177f
C11096 VDD.n3902 VSUBS 0.00299f
C11097 VDD.n3903 VSUBS 0.00134f
C11098 VDD.n3904 VSUBS 0.00627f
C11099 VDD.n3905 VSUBS 0.00194f
C11100 VDD.n3906 VSUBS 0.0155f
C11101 VDD.n3907 VSUBS 0.692f
C11102 VDD.n3908 VSUBS 0.0198f
C11103 VDD.n3909 VSUBS 0.539f
C11104 VDD.n3910 VSUBS 0.397f
C11105 VDD.n3911 VSUBS 0.0155f
C11106 VDD.n3912 VSUBS 0.173f
C11107 VDD.n3913 VSUBS 0.183f
C11108 VDD.n3914 VSUBS 0.00776f
C11109 VDD.n3915 VSUBS 0.00236f
C11110 VDD.n3916 VSUBS 0.00201f
C11111 VDD.n3917 VSUBS 0.00425f
C11112 VDD.n3918 VSUBS 0.00496f
C11113 VDD.n3919 VSUBS 0.00248f
C11114 VDD.n3920 VSUBS 0.00315f
C11115 VDD.n3921 VSUBS 0.00315f
C11116 VDD.n3922 VSUBS 0.00134f
C11117 VDD.n3923 VSUBS 0.0065f
C11118 VDD.n3924 VSUBS 0.00194f
C11119 VDD.t91 VSUBS 0.488f
C11120 VDD.n3925 VSUBS 0.0198f
C11121 VDD.n3926 VSUBS 0.163f
C11122 VDD.n3927 VSUBS 0.509f
C11123 VDD.n3928 VSUBS 0.0155f
C11124 VDD.n3929 VSUBS 0.173f
C11125 VDD.n3930 VSUBS 0.183f
C11126 VDD.n3931 VSUBS 0.00753f
C11127 VDD.n3932 VSUBS 0.00205f
C11128 VDD.n3933 VSUBS 0.00134f
C11129 VDD.n3934 VSUBS 5.9e-19
C11130 VDD.n3935 VSUBS 0.00153f
C11131 VDD.n3936 VSUBS 0.00248f
C11132 VDD.n3937 VSUBS 0.00401f
C11133 VDD.n3938 VSUBS 0.00507f
C11134 VDD.n3939 VSUBS 0.00224f
C11135 VDD.n3940 VSUBS 8.26e-19
C11136 VDD.n3941 VSUBS 0.0033f
C11137 VDD.n3942 VSUBS 0.0033f
C11138 VDD.n3943 VSUBS 0.00134f
C11139 VDD.n3944 VSUBS 0.00673f
C11140 VDD.n3945 VSUBS 0.00194f
C11141 VDD.n3946 VSUBS 0.0198f
C11142 VDD.n3947 VSUBS 0.539f
C11143 VDD.n3948 VSUBS 0.509f
C11144 VDD.n3949 VSUBS 0.0155f
C11145 VDD.n3950 VSUBS 0.173f
C11146 VDD.n3951 VSUBS 0.183f
C11147 VDD.n3952 VSUBS 0.0073f
C11148 VDD.n3953 VSUBS 0.00173f
C11149 VDD.n3954 VSUBS 0.00134f
C11150 VDD.n3955 VSUBS 0.00201f
C11151 VDD.n3956 VSUBS 0.00212f
C11152 VDD.n3957 VSUBS 0.00378f
C11153 VDD.n3958 VSUBS 0.0046f
C11154 VDD.n3959 VSUBS 0.00248f
C11155 VDD.n3960 VSUBS 0.00142f
C11156 VDD.n3961 VSUBS 0.00322f
C11157 VDD.n3962 VSUBS 0.00696f
C11158 VDD.n3963 VSUBS 0.00194f
C11159 VDD.n3964 VSUBS 0.0198f
C11160 VDD.n3965 VSUBS 0.539f
C11161 VDD.n3966 VSUBS 0.509f
C11162 VDD.n3967 VSUBS 0.0155f
C11163 VDD.n3968 VSUBS 0.153f
C11164 VDD.t11 VSUBS 0.0916f
C11165 VDD.n3969 VSUBS 0.112f
C11166 VDD.n3970 VSUBS 0.00707f
C11167 VDD.n3971 VSUBS 0.00134f
C11168 VDD.n3972 VSUBS 0.00134f
C11169 VDD.n3973 VSUBS 0.00201f
C11170 VDD.n3974 VSUBS 0.00201f
C11171 VDD.n3975 VSUBS 0.00346f
C11172 VDD.n3976 VSUBS 9.44e-19
C11173 VDD.n3977 VSUBS 7.08e-19
C11174 VDD.n3978 VSUBS 0.00354f
C11175 VDD.n3979 VSUBS 0.00413f
C11176 VDD.n3980 VSUBS 0.00271f
C11177 VDD.n3981 VSUBS 0.00189f
C11178 VDD.n3982 VSUBS 0.00307f
C11179 VDD.n3983 VSUBS 0.00134f
C11180 VDD.n3984 VSUBS 0.00201f
C11181 VDD.n3985 VSUBS 0.00189f
C11182 VDD.n3986 VSUBS 0.00106f
C11183 VDD.n3987 VSUBS 0.00719f
C11184 VDD.n3988 VSUBS 0.00194f
C11185 VDD.n3989 VSUBS 0.0198f
C11186 VDD.n3990 VSUBS 0.539f
C11187 VDD.n3991 VSUBS 0.509f
C11188 VDD.n3992 VSUBS 0.0155f
C11189 VDD.n3993 VSUBS 0.173f
C11190 VDD.n3994 VSUBS 0.183f
C11191 VDD.n3995 VSUBS 0.00684f
C11192 VDD.n3996 VSUBS 0.00126f
C11193 VDD.n3997 VSUBS 5.51e-19
C11194 VDD.n3998 VSUBS 5.51e-19
C11195 VDD.n3999 VSUBS 0.00346f
C11196 VDD.n4000 VSUBS 7.87e-19
C11197 VDD.n4001 VSUBS 0.00319f
C11198 VDD.n4002 VSUBS 0.00295f
C11199 VDD.n4003 VSUBS 0.00283f
C11200 VDD.n4004 VSUBS 0.00236f
C11201 VDD.n4005 VSUBS 0.00291f
C11202 VDD.n4006 VSUBS 0.00102f
C11203 VDD.n4007 VSUBS 0.00153f
C11204 VDD.n4008 VSUBS 0.00189f
C11205 VDD.n4009 VSUBS 0.0013f
C11206 VDD.n4010 VSUBS 0.00126f
C11207 VDD.n4011 VSUBS 0.00741f
C11208 VDD.n4012 VSUBS 0.00194f
C11209 VDD.n4013 VSUBS 0.0198f
C11210 VDD.n4014 VSUBS 0.539f
C11211 VDD.t72 VSUBS 0.387f
C11212 VDD.n4015 VSUBS 0.153f
C11213 VDD.n4016 VSUBS 0.0155f
C11214 VDD.n4017 VSUBS 0.173f
C11215 VDD.n4018 VSUBS 0.183f
C11216 VDD.n4019 VSUBS 0.00661f
C11217 VDD.n4020 VSUBS 7.08e-19
C11218 VDD.n4021 VSUBS 5.51e-19
C11219 VDD.n4022 VSUBS 0.00354f
C11220 VDD.n4023 VSUBS 9.44e-19
C11221 VDD.n4024 VSUBS 0.0033f
C11222 VDD.n4025 VSUBS 0.00283f
C11223 VDD.n4026 VSUBS 0.00283f
C11224 VDD.n4027 VSUBS 0.00134f
C11225 VDD.n4028 VSUBS 6.29e-19
C11226 VDD.n4029 VSUBS 0.00283f
C11227 VDD.n4030 VSUBS 0.0026f
C11228 VDD.n4031 VSUBS 9.44e-19
C11229 VDD.n4032 VSUBS 0.00201f
C11230 VDD.n4033 VSUBS 0.00177f
C11231 VDD.n4034 VSUBS 0.00764f
C11232 VDD.n4035 VSUBS 0.00194f
C11233 VDD.n4036 VSUBS 0.509f
C11234 VDD.n4037 VSUBS 0.509f
C11235 VDD.n4038 VSUBS 0.0155f
C11236 VDD.n4039 VSUBS 0.173f
C11237 VDD.n4040 VSUBS 0.183f
C11238 VDD.n4041 VSUBS 0.00639f
C11239 VDD.n4042 VSUBS 0.00102f
C11240 VDD.n4043 VSUBS 3.93e-19
C11241 VDD.n4044 VSUBS 0.00378f
C11242 VDD.n4045 VSUBS 0.0011f
C11243 VDD.n4046 VSUBS 0.0026f
C11244 VDD.n4047 VSUBS 0.00307f
C11245 VDD.n4048 VSUBS 0.00366f
C11246 VDD.n4049 VSUBS 0.00307f
C11247 VDD.n4050 VSUBS 0.00295f
C11248 VDD.n4051 VSUBS 0.00134f
C11249 VDD.n4052 VSUBS 0.00201f
C11250 VDD.n4053 VSUBS 0.00201f
C11251 VDD.n4054 VSUBS 0.00593f
C11252 VDD.n4055 VSUBS 0.00194f
C11253 VDD.n4056 VSUBS 0.539f
C11254 VDD.n4057 VSUBS 0.377f
C11255 VDD.n4058 VSUBS 0.173f
C11256 VDD.n4059 VSUBS 0.183f
C11257 VDD.n4060 VSUBS 0.00616f
C11258 VDD.n4061 VSUBS 0.00118f
C11259 VDD.n4062 VSUBS 2.36e-19
C11260 VDD.n4063 VSUBS 0.00393f
C11261 VDD.n4064 VSUBS 0.00126f
C11262 VDD.n4065 VSUBS 0.00189f
C11263 VDD.n4066 VSUBS 0.00307f
C11264 VDD.n4067 VSUBS 0.00637f
C11265 VDD.n4068 VSUBS 0.00496f
C11266 VDD.n4069 VSUBS 0.00409f
C11267 VDD.n4070 VSUBS 0.00134f
C11268 VDD.n4071 VSUBS 0.00593f
C11269 VDD.n4072 VSUBS 0.00194f
C11270 VDD.t47 VSUBS 0.346f
C11271 VDD.n4073 VSUBS 0.153f
C11272 VDD.n4074 VSUBS 0.183f
C11273 VDD.n4075 VSUBS 0.173f
C11274 VDD.n4076 VSUBS 0.509f
C11275 VDD.n4077 VSUBS 0.00616f
C11276 VDD.n4078 VSUBS 1.57e-19
C11277 VDD.n4079 VSUBS 0.00134f
C11278 VDD.n4080 VSUBS 0.00118f
C11279 VDD.n4081 VSUBS 0.00189f
C11280 VDD.n4082 VSUBS 0.00409f
C11281 VDD.n4083 VSUBS 0.00201f
C11282 VDD.n4084 VSUBS 0.00413f
C11283 VDD.n4085 VSUBS 0.00507f
C11284 VDD.n4086 VSUBS 0.00248f
C11285 VDD.n4087 VSUBS 0.00393f
C11286 VDD.n4088 VSUBS 0.00134f
C11287 VDD.n4089 VSUBS 0.00764f
C11288 VDD.n4090 VSUBS 0.00194f
C11289 VDD.n4091 VSUBS 0.539f
C11290 VDD.n4092 VSUBS 0.183f
C11291 VDD.n4093 VSUBS 0.173f
C11292 VDD.n4094 VSUBS 0.509f
C11293 VDD.n4095 VSUBS 0.00639f
C11294 VDD.n4096 VSUBS 4.72e-19
C11295 VDD.n4097 VSUBS 0.00393f
C11296 VDD.n4098 VSUBS 0.00134f
C11297 VDD.n4099 VSUBS 4.72e-19
C11298 VDD.n4100 VSUBS 0.00165f
C11299 VDD.n4101 VSUBS 0.00248f
C11300 VDD.n4102 VSUBS 0.00389f
C11301 VDD.n4103 VSUBS 0.00507f
C11302 VDD.n4104 VSUBS 0.00236f
C11303 VDD.n4105 VSUBS 8.26e-19
C11304 VDD.n4106 VSUBS 0.00378f
C11305 VDD.n4107 VSUBS 0.00134f
C11306 VDD.n4108 VSUBS 0.00741f
C11307 VDD.n4109 VSUBS 0.00194f
C11308 VDD.n4110 VSUBS 0.539f
C11309 VDD.n4111 VSUBS 0.0916f
C11310 VDD.t135 VSUBS 0.122f
C11311 VDD.n4112 VSUBS 0.142f
C11312 VDD.n4113 VSUBS 0.509f
C11313 VDD.n4114 VSUBS 0.00661f
C11314 VDD.n4115 VSUBS 7.87e-19
C11315 VDD.n4116 VSUBS 0.00378f
C11316 VDD.n4117 VSUBS 0.00134f
C11317 VDD.n4118 VSUBS 0.00201f
C11318 VDD.n4119 VSUBS 0.00212f
C11319 VDD.n4120 VSUBS 0.00366f
C11320 VDD.n4121 VSUBS 0.0046f
C11321 VDD.n4122 VSUBS 0.0026f
C11322 VDD.n4123 VSUBS 0.00142f
C11323 VDD.n4124 VSUBS 0.00362f
C11324 VDD.n4125 VSUBS 0.00134f
C11325 VDD.n4126 VSUBS 0.00719f
C11326 VDD.n4127 VSUBS 0.00194f
C11327 VDD.n4128 VSUBS 0.539f
C11328 VDD.n4129 VSUBS 0.183f
C11329 VDD.n4130 VSUBS 0.173f
C11330 VDD.n4131 VSUBS 0.509f
C11331 VDD.n4132 VSUBS 0.00684f
C11332 VDD.n4133 VSUBS 8.65e-19
C11333 VDD.n4134 VSUBS 0.00134f
C11334 VDD.n4135 VSUBS 0.00134f
C11335 VDD.n4136 VSUBS 0.00201f
C11336 VDD.n4137 VSUBS 0.00201f
C11337 VDD.n4138 VSUBS 0.00283f
C11338 VDD.n4139 VSUBS 0.00342f
C11339 VDD.n4140 VSUBS 0.00413f
C11340 VDD.n4141 VSUBS 0.00283f
C11341 VDD.n4142 VSUBS 0.00189f
C11342 VDD.n4143 VSUBS 0.00315f
C11343 VDD.n4144 VSUBS 0.00134f
C11344 VDD.n4145 VSUBS 0.00696f
C11345 VDD.n4146 VSUBS 0.00194f
C11346 VDD.n4147 VSUBS 0.539f
C11347 VDD.n4148 VSUBS 0.183f
C11348 VDD.n4149 VSUBS 0.173f
C11349 VDD.t133 VSUBS 0.417f
C11350 VDD.n4150 VSUBS 0.132f
C11351 VDD.n4151 VSUBS 0.00707f
C11352 VDD.n4152 VSUBS 8.65e-19
C11353 VDD.n4153 VSUBS 0.00134f
C11354 VDD.n4154 VSUBS 0.00201f
C11355 VDD.n4155 VSUBS 0.00189f
C11356 VDD.n4156 VSUBS 9.44e-19
C11357 VDD.n4157 VSUBS 0.00126f
C11358 VDD.n4158 VSUBS 6.29e-19
C11359 VDD.n4159 VSUBS 0.00275f
C11360 VDD.n4160 VSUBS 0.00319f
C11361 VDD.n4161 VSUBS 0.00295f
C11362 VDD.n4162 VSUBS 0.00295f
C11363 VDD.n4163 VSUBS 0.00267f
C11364 VDD.n4164 VSUBS 0.00134f
C11365 VDD.n4165 VSUBS 0.00134f
C11366 VDD.n4166 VSUBS 0.00673f
C11367 VDD.n4167 VSUBS 0.00194f
C11368 VDD.n4168 VSUBS 0.499f
C11369 VDD.n4169 VSUBS 0.183f
C11370 VDD.n4170 VSUBS 0.173f
C11371 VDD.n4171 VSUBS 0.539f
C11372 VDD.n4172 VSUBS 0.509f
C11373 VDD.n4173 VSUBS 0.0073f
C11374 VDD.n4174 VSUBS 0.00181f
C11375 VDD.n4175 VSUBS 0.00378f
C11376 VDD.n4176 VSUBS 0.00201f
C11377 VDD.n4177 VSUBS 0.0013f
C11378 VDD.n4178 VSUBS 8.65e-19
C11379 VDD.n4179 VSUBS 0.00283f
C11380 VDD.n4180 VSUBS 0.00319f
C11381 VDD.n4181 VSUBS 0.00283f
C11382 VDD.n4182 VSUBS 0.00283f
C11383 VDD.n4183 VSUBS 0.00267f
C11384 VDD.n4184 VSUBS 0.00118f
C11385 VDD.n4185 VSUBS 0.00134f
C11386 VDD.n4186 VSUBS 0.0065f
C11387 VDD.n4187 VSUBS 0.00194f
C11388 VDD.n4188 VSUBS 0.183f
C11389 VDD.n4189 VSUBS 0.173f
C11390 VDD.n4190 VSUBS 0.315f
C11391 VDD.t33 VSUBS 0.377f
C11392 VDD.n4191 VSUBS 0.356f
C11393 VDD.n4192 VSUBS 0.00753f
C11394 VDD.n4193 VSUBS 6.29e-19
C11395 VDD.n4194 VSUBS 0.00102f
C11396 VDD.n4195 VSUBS 0.00271f
C11397 VDD.n4196 VSUBS 9.44e-19
C11398 VDD.n4197 VSUBS 0.00201f
C11399 VDD.n4198 VSUBS 0.00177f
C11400 VDD.n4199 VSUBS 0.00118f
C11401 VDD.n4200 VSUBS 0.00283f
C11402 VDD.n4201 VSUBS 0.00248f
C11403 VDD.n4202 VSUBS 0.00307f
C11404 VDD.n4203 VSUBS 0.00378f
C11405 VDD.n4204 VSUBS 0.00267f
C11406 VDD.n4205 VSUBS 0.00134f
C11407 VDD.n4206 VSUBS 0.00627f
C11408 VDD.n4207 VSUBS 0.00194f
C11409 VDD.n4208 VSUBS 0.183f
C11410 VDD.n4209 VSUBS 0.173f
C11411 VDD.n4210 VSUBS 0.692f
C11412 VDD.n4211 VSUBS 0.539f
C11413 VDD.n4212 VSUBS 0.509f
C11414 VDD.n4213 VSUBS 0.00776f
C11415 VDD.n4214 VSUBS 0.00134f
C11416 VDD.n4215 VSUBS 0.00295f
C11417 VDD.n4216 VSUBS 0.00134f
C11418 VDD.n4217 VSUBS 0.00201f
C11419 VDD.n4218 VSUBS 0.00201f
C11420 VDD.n4219 VSUBS 0.00134f
C11421 VDD.n4220 VSUBS 0.00283f
C11422 VDD.n4221 VSUBS 0.00177f
C11423 VDD.n4222 VSUBS 0.00307f
C11424 VDD.n4223 VSUBS 0.00649f
C11425 VDD.n4224 VSUBS 0.0138f
C11426 VDD.n4225 VSUBS 0.00535f
C11427 VDD.n4226 VSUBS 0.0138f
C11428 VDD.n4227 VSUBS 0.00551f
C11429 VDD.n4228 VSUBS 0.00535f
C11430 VDD.n4229 VSUBS 0.00602f
C11431 VDD.n4230 VSUBS 0.00307f
C11432 VDD.n4231 VSUBS 0.00496f
C11433 VDD.n4232 VSUBS 0.00519f
C11434 VDD.n4233 VSUBS 0.00248f
C11435 VDD.n4234 VSUBS 0.00299f
C11436 VDD.n4235 VSUBS 0.00134f
C11437 VDD.n4236 VSUBS 3.54e-19
C11438 VDD.n4237 VSUBS 0.00177f
C11439 VDD.n4238 VSUBS 0.00299f
C11440 VDD.n4239 VSUBS 0.00134f
C11441 VDD.n4240 VSUBS 0.00627f
C11442 VDD.n4241 VSUBS 0.00194f
C11443 VDD.n4242 VSUBS 0.58f
C11444 VDD.t105 VSUBS 0.183f
C11445 VDD.n4243 VSUBS 0.621f
C11446 VDD.n4244 VSUBS 0.539f
C11447 VDD.n4245 VSUBS 0.509f
C11448 VDD.n4246 VSUBS 0.173f
C11449 VDD.n4247 VSUBS 0.183f
C11450 VDD.n4248 VSUBS 0.00776f
C11451 VDD.n4249 VSUBS 0.00236f
C11452 VDD.n4250 VSUBS 0.00248f
C11453 VDD.n4251 VSUBS 0.00378f
C11454 VDD.n4252 VSUBS 0.00507f
C11455 VDD.n4253 VSUBS 0.00248f
C11456 VDD.n4254 VSUBS 8.26e-19
C11457 VDD.n4255 VSUBS 0.00315f
C11458 VDD.n4256 VSUBS 0.00315f
C11459 VDD.n4257 VSUBS 0.00134f
C11460 VDD.n4258 VSUBS 0.0065f
C11461 VDD.n4259 VSUBS 0.00194f
C11462 VDD.n4260 VSUBS 0.539f
C11463 VDD.t13 VSUBS 0.468f
C11464 VDD.n4261 VSUBS 0.112f
C11465 VDD.n4262 VSUBS 0.173f
C11466 VDD.n4263 VSUBS 0.183f
C11467 VDD.n4264 VSUBS 0.00753f
C11468 VDD.n4265 VSUBS 0.00205f
C11469 VDD.n4266 VSUBS 0.00134f
C11470 VDD.n4267 VSUBS 0.00201f
C11471 VDD.n4268 VSUBS 0.00212f
C11472 VDD.n4269 VSUBS 0.00354f
C11473 VDD.n4270 VSUBS 0.0046f
C11474 VDD.n4271 VSUBS 0.00271f
C11475 VDD.n4272 VSUBS 0.00142f
C11476 VDD.n4273 VSUBS 0.00307f
C11477 VDD.n4274 VSUBS 0.00673f
C11478 VDD.n4275 VSUBS 0.00194f
C11479 VDD.n4276 VSUBS 0.468f
C11480 VDD.n4277 VSUBS 0.509f
C11481 VDD.n4278 VSUBS 0.173f
C11482 VDD.n4279 VSUBS 0.183f
C11483 VDD.n4280 VSUBS 0.0073f
C11484 VDD.n4281 VSUBS 0.00134f
C11485 VDD.n4282 VSUBS 0.00134f
C11486 VDD.n4283 VSUBS 0.00201f
C11487 VDD.n4284 VSUBS 0.00201f
C11488 VDD.n4285 VSUBS 0.0033f
C11489 VDD.n4286 VSUBS 0.0011f
C11490 VDD.n4287 VSUBS 8.65e-19
C11491 VDD.n4288 VSUBS 0.0033f
C11492 VDD.n4289 VSUBS 0.00413f
C11493 VDD.n4290 VSUBS 0.00295f
C11494 VDD.n4291 VSUBS 0.00189f
C11495 VDD.n4292 VSUBS 0.00291f
C11496 VDD.n4293 VSUBS 0.00134f
C11497 VDD.n4294 VSUBS 0.00201f
C11498 VDD.n4295 VSUBS 0.00696f
C11499 VDD.n4296 VSUBS 0.00194f
C11500 VDD.n4297 VSUBS 0.539f
C11501 VDD.n4298 VSUBS 0.336f
C11502 VDD.n4299 VSUBS 0.173f
C11503 VDD.n4300 VSUBS 0.183f
C11504 VDD.n4301 VSUBS 0.00707f
C11505 VDD.n4302 VSUBS 0.00181f
C11506 VDD.n4303 VSUBS 0.00271f
C11507 VDD.n4304 VSUBS 0.00338f
C11508 VDD.n4305 VSUBS 7.87e-19
C11509 VDD.n4306 VSUBS 7.08e-19
C11510 VDD.n4307 VSUBS 0.00319f
C11511 VDD.n4308 VSUBS 0.00295f
C11512 VDD.n4309 VSUBS 0.00295f
C11513 VDD.n4310 VSUBS 9.44e-19
C11514 VDD.n4311 VSUBS 0.00283f
C11515 VDD.n4312 VSUBS 0.00248f
C11516 VDD.n4313 VSUBS 0.00142f
C11517 VDD.n4314 VSUBS 0.00201f
C11518 VDD.n4315 VSUBS 0.0013f
C11519 VDD.n4316 VSUBS 0.00134f
C11520 VDD.n4317 VSUBS 0.00719f
C11521 VDD.n4318 VSUBS 0.00194f
C11522 VDD.t129 VSUBS 0.427f
C11523 VDD.n4319 VSUBS 0.285f
C11524 VDD.n4320 VSUBS 0.509f
C11525 VDD.n4321 VSUBS 0.173f
C11526 VDD.n4322 VSUBS 0.183f
C11527 VDD.n4323 VSUBS 0.00684f
C11528 VDD.n4324 VSUBS 8.65e-19
C11529 VDD.n4325 VSUBS 0.00338f
C11530 VDD.n4326 VSUBS 9.44e-19
C11531 VDD.n4327 VSUBS 5.51e-19
C11532 VDD.n4328 VSUBS 0.00307f
C11533 VDD.n4329 VSUBS 0.00283f
C11534 VDD.n4330 VSUBS 0.00283f
C11535 VDD.n4331 VSUBS 0.00134f
C11536 VDD.n4332 VSUBS 6.29e-19
C11537 VDD.n4333 VSUBS 0.00283f
C11538 VDD.n4334 VSUBS 0.00283f
C11539 VDD.n4335 VSUBS 9.44e-19
C11540 VDD.n4336 VSUBS 0.00201f
C11541 VDD.n4337 VSUBS 0.00177f
C11542 VDD.n4338 VSUBS 0.00741f
C11543 VDD.n4339 VSUBS 0.00194f
C11544 VDD.n4340 VSUBS 0.539f
C11545 VDD.n4341 VSUBS 0.509f
C11546 VDD.n4342 VSUBS 0.173f
C11547 VDD.n4343 VSUBS 0.183f
C11548 VDD.n4344 VSUBS 0.00661f
C11549 VDD.n4345 VSUBS 0.00118f
C11550 VDD.n4346 VSUBS 0.00378f
C11551 VDD.n4347 VSUBS 0.0011f
C11552 VDD.n4348 VSUBS 3.93e-19
C11553 VDD.n4349 VSUBS 0.00236f
C11554 VDD.n4350 VSUBS 0.00307f
C11555 VDD.n4351 VSUBS 0.00389f
C11556 VDD.n4352 VSUBS 0.00291f
C11557 VDD.n4353 VSUBS 0.00295f
C11558 VDD.n4354 VSUBS 0.00134f
C11559 VDD.n4355 VSUBS 0.00201f
C11560 VDD.n4356 VSUBS 0.00201f
C11561 VDD.n4357 VSUBS 0.00764f
C11562 VDD.n4358 VSUBS 0.00194f
C11563 VDD.n4359 VSUBS 0.438f
C11564 VDD.t78 VSUBS 0.153f
C11565 VDD.n4360 VSUBS 0.509f
C11566 VDD.n4361 VSUBS 0.173f
C11567 VDD.n4362 VSUBS 0.132f
C11568 VDD.n4363 VSUBS 0.00639f
C11569 VDD.n4364 VSUBS 0.00134f
C11570 VDD.n4365 VSUBS 0.00393f
C11571 VDD.n4366 VSUBS 0.00126f
C11572 VDD.n4367 VSUBS 2.36e-19
C11573 VDD.n4368 VSUBS 0.00165f
C11574 VDD.n4369 VSUBS 0.00307f
C11575 VDD.n4370 VSUBS 0.0046f
C11576 VDD.n4371 VSUBS 0.00409f
C11577 VDD.n4372 VSUBS 0.00496f
C11578 VDD.n4373 VSUBS 0.00409f
C11579 VDD.n4374 VSUBS 0.00134f
C11580 VDD.n4375 VSUBS 0.00593f
C11581 VDD.n4376 VSUBS 0.00194f
C11582 VDD.n4377 VSUBS 0.539f
C11583 VDD.n4378 VSUBS 0.509f
C11584 VDD.n4379 VSUBS 0.173f
C11585 VDD.n4380 VSUBS 0.183f
C11586 VDD.n4381 VSUBS 0.00616f
C11587 VDD.n4382 VSUBS 1.57e-19
C11588 VDD.n4383 VSUBS 0.00134f
C11589 VDD.n4384 VSUBS 0.00201f
C11590 VDD.n4385 VSUBS 0.00106f
C11591 VDD.n4386 VSUBS 0.00295f
C11592 VDD.n4387 VSUBS 0.00496f
C11593 VDD.n4388 VSUBS 0.00531f
C11594 VDD.n4389 VSUBS 0.00248f
C11595 VDD.n4390 VSUBS 0.00409f
C11596 VDD.n4391 VSUBS 0.00134f
C11597 VDD.n4392 VSUBS 0.00593f
C11598 VDD.n4393 VSUBS 0.00194f
C11599 VDD.n4394 VSUBS 0.366f
C11600 VDD.n4395 VSUBS 0.183f
C11601 VDD.n4396 VSUBS 0.173f
C11602 VDD.t27 VSUBS 0.499f
C11603 VDD.n4397 VSUBS 0.0916f
C11604 VDD.n4398 VSUBS 0.00616f
C11605 VDD.n4399 VSUBS 1.57e-19
C11606 VDD.n4400 VSUBS 0.00134f
C11607 VDD.n4401 VSUBS 2.36e-19
C11608 VDD.n4402 VSUBS 0.00189f
C11609 VDD.n4403 VSUBS 0.00409f
C11610 VDD.n4404 VSUBS 0.00248f
C11611 VDD.n4405 VSUBS 0.00366f
C11612 VDD.n4406 VSUBS 0.00507f
C11613 VDD.n4407 VSUBS 0.0026f
C11614 VDD.n4408 VSUBS 8.26e-19
C11615 VDD.n4409 VSUBS 0.00393f
C11616 VDD.n4410 VSUBS 0.00134f
C11617 VDD.n4411 VSUBS 0.00764f
C11618 VDD.n4412 VSUBS 0.00194f
C11619 VDD.n4413 VSUBS 0.458f
C11620 VDD.n4414 VSUBS 0.183f
C11621 VDD.n4415 VSUBS 0.173f
C11622 VDD.n4416 VSUBS 0.509f
C11623 VDD.n4417 VSUBS 0.00639f
C11624 VDD.n4418 VSUBS 4.72e-19
C11625 VDD.n4419 VSUBS 0.00393f
C11626 VDD.n4420 VSUBS 0.00134f
C11627 VDD.n4421 VSUBS 0.00201f
C11628 VDD.n4422 VSUBS 0.00212f
C11629 VDD.n4423 VSUBS 0.00342f
C11630 VDD.n4424 VSUBS 0.0046f
C11631 VDD.n4425 VSUBS 0.00283f
C11632 VDD.n4426 VSUBS 0.00142f
C11633 VDD.n4427 VSUBS 0.00378f
C11634 VDD.n4428 VSUBS 0.00134f
C11635 VDD.n4429 VSUBS 0.00741f
C11636 VDD.n4430 VSUBS 0.00194f
C11637 VDD.n4431 VSUBS 0.539f
C11638 VDD.n4432 VSUBS 0.183f
C11639 VDD.n4433 VSUBS 0.173f
C11640 VDD.t70 VSUBS 0.458f
C11641 VDD.n4434 VSUBS 0.315f
C11642 VDD.n4435 VSUBS 0.00661f
C11643 VDD.n4436 VSUBS 5.51e-19
C11644 VDD.n4437 VSUBS 0.00134f
C11645 VDD.n4438 VSUBS 0.00201f
C11646 VDD.n4439 VSUBS 0.00134f
C11647 VDD.n4440 VSUBS 0.00201f
C11648 VDD.n4441 VSUBS 0.00283f
C11649 VDD.n4442 VSUBS 0.00319f
C11650 VDD.n4443 VSUBS 0.00413f
C11651 VDD.n4444 VSUBS 0.00307f
C11652 VDD.n4445 VSUBS 0.00346f
C11653 VDD.n4446 VSUBS 0.00134f
C11654 VDD.n4447 VSUBS 0.00719f
C11655 VDD.n4448 VSUBS 0.00194f
C11656 VDD.n4449 VSUBS 0.275f
C11657 VDD.n4450 VSUBS 0.183f
C11658 VDD.n4451 VSUBS 0.0155f
C11659 VDD.n4452 VSUBS 0.173f
C11660 VDD.n4453 VSUBS 0.509f
C11661 VDD.n4454 VSUBS 0.00684f
C11662 VDD.n4455 VSUBS 0.00181f
C11663 VDD.n4456 VSUBS 0.00378f
C11664 VDD.n4457 VSUBS 0.00201f
C11665 VDD.n4458 VSUBS 8.26e-19
C11666 VDD.n4459 VSUBS 0.00134f
C11667 VDD.n4460 VSUBS 5.51e-19
C11668 VDD.n4461 VSUBS 0.00283f
C11669 VDD.n4462 VSUBS 0.00307f
C11670 VDD.n4463 VSUBS 0.00295f
C11671 VDD.n4464 VSUBS 0.00295f
C11672 VDD.n4465 VSUBS 0.00299f
C11673 VDD.n4466 VSUBS 0.00118f
C11674 VDD.n4467 VSUBS 0.00696f
C11675 VDD.n4468 VSUBS 0.00194f
C11676 VDD.n4469 VSUBS 0.0198f
C11677 VDD.n4470 VSUBS 0.539f
C11678 VDD.n4471 VSUBS 0.183f
C11679 VDD.n4472 VSUBS 0.0155f
C11680 VDD.n4473 VSUBS 0.173f
C11681 VDD.n4474 VSUBS 0.509f
C11682 VDD.n4475 VSUBS 0.00707f
C11683 VDD.n4476 VSUBS 9.44e-19
C11684 VDD.n4477 VSUBS 7.08e-19
C11685 VDD.n4478 VSUBS 0.0026f
C11686 VDD.n4479 VSUBS 0.00142f
C11687 VDD.n4480 VSUBS 0.00201f
C11688 VDD.n4481 VSUBS 0.0013f
C11689 VDD.n4482 VSUBS 0.00134f
C11690 VDD.n4483 VSUBS 8.65e-19
C11691 VDD.n4484 VSUBS 0.00283f
C11692 VDD.n4485 VSUBS 0.00295f
C11693 VDD.n4486 VSUBS 0.00283f
C11694 VDD.n4487 VSUBS 0.00283f
C11695 VDD.n4488 VSUBS 0.00299f
C11696 VDD.n4489 VSUBS 0.00102f
C11697 VDD.n4490 VSUBS 0.00134f
C11698 VDD.n4491 VSUBS 0.00673f
C11699 VDD.n4492 VSUBS 0.00194f
C11700 VDD.n4493 VSUBS 0.0198f
C11701 VDD.n4494 VSUBS 0.448f
C11702 VDD.t110 VSUBS 0.122f
C11703 VDD.n4495 VSUBS 0.153f
C11704 VDD.n4496 VSUBS 0.0155f
C11705 VDD.n4497 VSUBS 0.173f
C11706 VDD.n4498 VSUBS 0.509f
C11707 VDD.n4499 VSUBS 0.0073f
C11708 VDD.n4500 VSUBS 6.29e-19
C11709 VDD.n4501 VSUBS 8.65e-19
C11710 VDD.n4502 VSUBS 0.00295f
C11711 VDD.n4503 VSUBS 9.44e-19
C11712 VDD.n4504 VSUBS 0.00201f
C11713 VDD.n4505 VSUBS 0.00177f
C11714 VDD.n4506 VSUBS 0.00118f
C11715 VDD.n4507 VSUBS 0.00283f
C11716 VDD.n4508 VSUBS 0.00224f
C11717 VDD.n4509 VSUBS 0.00307f
C11718 VDD.n4510 VSUBS 0.00401f
C11719 VDD.n4511 VSUBS 0.00299f
C11720 VDD.n4512 VSUBS 0.00134f
C11721 VDD.n4513 VSUBS 0.0065f
C11722 VDD.n4514 VSUBS 0.00194f
C11723 VDD.n4515 VSUBS 0.0198f
C11724 VDD.n4516 VSUBS 0.539f
C11725 VDD.n4517 VSUBS 0.183f
C11726 VDD.n4518 VSUBS 0.0155f
C11727 VDD.n4519 VSUBS 0.173f
C11728 VDD.n4520 VSUBS 0.0198f
C11729 VDD.n4521 VSUBS 0.539f
C11730 VDD.n4522 VSUBS 0.509f
C11731 VDD.n4523 VSUBS 0.00753f
C11732 VDD.n4524 VSUBS 0.00236f
C11733 VDD.n4525 VSUBS 0.00496f
C11734 VDD.n4526 VSUBS 0.00299f
C11735 VDD.n4527 VSUBS 0.00417f
C11736 VDD.n4528 VSUBS 0.00354f
C11737 VDD.n4529 VSUBS 0.00307f
C11738 VDD.n4530 VSUBS 0.00472f
C11739 VDD.n4531 VSUBS 0.00496f
C11740 VDD.n4532 VSUBS 0.00134f
C11741 VDD.n4533 VSUBS 0.00627f
C11742 VDD.n4534 VSUBS 0.00194f
C11743 VDD.n4535 VSUBS 0.183f
C11744 VDD.n4536 VSUBS 0.0155f
C11745 VDD.n4537 VSUBS 0.0916f
C11746 VDD.t50 VSUBS 0.153f
C11747 VDD.n4538 VSUBS 0.0155f
C11748 VDD.n4539 VSUBS 0.692f
C11749 VDD.n4540 VSUBS 0.0198f
C11750 VDD.n4541 VSUBS 0.539f
C11751 VDD.n4542 VSUBS 0.438f
C11752 VDD.n4543 VSUBS 0.00776f
C11753 VDD.n4544 VSUBS 0.00236f
C11754 VDD.n4545 VSUBS 0.00299f
C11755 VDD.n4546 VSUBS 0.00134f
C11756 VDD.n4547 VSUBS 0.00201f
C11757 VDD.n4548 VSUBS 0.00106f
C11758 VDD.n4549 VSUBS 0.00283f
C11759 VDD.n4550 VSUBS 0.00496f
C11760 VDD.n4551 VSUBS 0.00543f
C11761 VDD.n4552 VSUBS 0.0138f
C11762 VDD.n4553 VSUBS 0.00551f
C11763 VDD.n4554 VSUBS 0.0138f
C11764 VDD.n4555 VSUBS 0.00551f
C11765 VDD.n4556 VSUBS 0.00535f
C11766 VDD.n4557 VSUBS 0.0026f
C11767 VDD.n4558 VSUBS 0.0026f
C11768 VDD.n4559 VSUBS 0.00543f
C11769 VDD.n4560 VSUBS 0.00507f
C11770 VDD.n4561 VSUBS 0.00271f
C11771 VDD.n4562 VSUBS 8.26e-19
C11772 VDD.n4563 VSUBS 0.00299f
C11773 VDD.n4564 VSUBS 0.00134f
C11774 VDD.n4565 VSUBS 0.00201f
C11775 VDD.n4566 VSUBS 0.00299f
C11776 VDD.n4567 VSUBS 0.00134f
C11777 VDD.n4568 VSUBS 0.00627f
C11778 VDD.n4569 VSUBS 0.00194f
C11779 VDD.n4570 VSUBS 0.0198f
C11780 VDD.n4571 VSUBS 0.692f
C11781 VDD.n4572 VSUBS 0.0155f
C11782 VDD.n4573 VSUBS 0.478f
C11783 VDD.t21 VSUBS 0.509f
C11784 VDD.n4574 VSUBS 0.0198f
C11785 VDD.n4575 VSUBS 0.244f
C11786 VDD.n4576 VSUBS 0.509f
C11787 VDD.n4577 VSUBS 0.0155f
C11788 VDD.n4578 VSUBS 0.173f
C11789 VDD.n4579 VSUBS 0.183f
C11790 VDD.n4580 VSUBS 0.00776f
C11791 VDD.n4581 VSUBS 0.00236f
C11792 VDD.n4582 VSUBS 0.00212f
C11793 VDD.n4583 VSUBS 0.0033f
C11794 VDD.n4584 VSUBS 0.0046f
C11795 VDD.n4585 VSUBS 0.00295f
C11796 VDD.n4586 VSUBS 0.00142f
C11797 VDD.n4587 VSUBS 0.00291f
C11798 VDD.n4588 VSUBS 0.00134f
C11799 VDD.n4589 VSUBS 0.00201f
C11800 VDD.n4590 VSUBS 0.0065f
C11801 VDD.n4591 VSUBS 0.00194f
C11802 VDD.n4592 VSUBS 0.0198f
C11803 VDD.n4593 VSUBS 0.539f
C11804 VDD.n4594 VSUBS 0.509f
C11805 VDD.n4595 VSUBS 0.0155f
C11806 VDD.n4596 VSUBS 0.173f
C11807 VDD.n4597 VSUBS 0.183f
C11808 VDD.n4598 VSUBS 0.00753f
C11809 VDD.n4599 VSUBS 0.00134f
C11810 VDD.n4600 VSUBS 0.00201f
C11811 VDD.n4601 VSUBS 0.00307f
C11812 VDD.n4602 VSUBS 0.00126f
C11813 VDD.n4603 VSUBS 0.00102f
C11814 VDD.n4604 VSUBS 0.00307f
C11815 VDD.n4605 VSUBS 0.00413f
C11816 VDD.n4606 VSUBS 0.00307f
C11817 VDD.n4607 VSUBS 0.00126f
C11818 VDD.n4608 VSUBS 0.00283f
C11819 VDD.n4609 VSUBS 0.00201f
C11820 VDD.n4610 VSUBS 0.00189f
C11821 VDD.n4611 VSUBS 0.00201f
C11822 VDD.n4612 VSUBS 8.26e-19
C11823 VDD.n4613 VSUBS 0.00134f
C11824 VDD.n4614 VSUBS 0.00673f
C11825 VDD.n4615 VSUBS 0.00194f
C11826 VDD.n4616 VSUBS 0.0198f
C11827 VDD.n4617 VSUBS 0.478f
C11828 VDD.t115 VSUBS 0.0712f
C11829 VDD.n4618 VSUBS 0.509f
C11830 VDD.n4619 VSUBS 0.0155f
C11831 VDD.n4620 VSUBS 0.173f
C11832 VDD.n4621 VSUBS 0.173f
C11833 VDD.n4622 VSUBS 0.0073f
C11834 VDD.n4623 VSUBS 5.51e-19
C11835 VDD.n4624 VSUBS 0.00307f
C11836 VDD.n4625 VSUBS 9.44e-19
C11837 VDD.n4626 VSUBS 8.65e-19
C11838 VDD.n4627 VSUBS 0.00295f
C11839 VDD.n4628 VSUBS 0.00295f
C11840 VDD.n4629 VSUBS 0.00295f
C11841 VDD.n4630 VSUBS 9.44e-19
C11842 VDD.n4631 VSUBS 0.00283f
C11843 VDD.n4632 VSUBS 0.00271f
C11844 VDD.n4633 VSUBS 0.00142f
C11845 VDD.n4634 VSUBS 0.00201f
C11846 VDD.n4635 VSUBS 0.0013f
C11847 VDD.n4636 VSUBS 0.00134f
C11848 VDD.n4637 VSUBS 0.00696f
C11849 VDD.n4638 VSUBS 0.00194f
C11850 VDD.n4639 VSUBS 0.0198f
C11851 VDD.n4640 VSUBS 0.539f
C11852 VDD.n4641 VSUBS 0.509f
C11853 VDD.n4642 VSUBS 0.0155f
C11854 VDD.n4643 VSUBS 0.173f
C11855 VDD.n4644 VSUBS 0.183f
C11856 VDD.n4645 VSUBS 0.00707f
C11857 VDD.n4646 VSUBS 8.65e-19
C11858 VDD.n4647 VSUBS 0.00307f
C11859 VDD.n4648 VSUBS 0.0011f
C11860 VDD.n4649 VSUBS 7.08e-19
C11861 VDD.n4650 VSUBS 0.00283f
C11862 VDD.n4651 VSUBS 0.00283f
C11863 VDD.n4652 VSUBS 0.00283f
C11864 VDD.n4653 VSUBS 0.00134f
C11865 VDD.n4654 VSUBS 6.29e-19
C11866 VDD.n4655 VSUBS 0.00283f
C11867 VDD.n4656 VSUBS 0.00307f
C11868 VDD.n4657 VSUBS 9.44e-19
C11869 VDD.n4658 VSUBS 0.00201f
C11870 VDD.n4659 VSUBS 0.00177f
C11871 VDD.n4660 VSUBS 0.00719f
C11872 VDD.n4661 VSUBS 0.00194f
C11873 VDD.n4662 VSUBS 0.0198f
C11874 VDD.n4663 VSUBS 0.539f
C11875 VDD.n4664 VSUBS 0.458f
C11876 VDD.t93 VSUBS 0.102f
C11877 VDD.n4665 VSUBS 0.0155f
C11878 VDD.n4666 VSUBS 0.122f
C11879 VDD.n4667 VSUBS 0.183f
C11880 VDD.n4668 VSUBS 0.00684f
C11881 VDD.n4669 VSUBS 0.00118f
C11882 VDD.n4670 VSUBS 0.00354f
C11883 VDD.n4671 VSUBS 0.00126f
C11884 VDD.n4672 VSUBS 5.51e-19
C11885 VDD.n4673 VSUBS 0.00212f
C11886 VDD.n4674 VSUBS 0.00307f
C11887 VDD.n4675 VSUBS 0.00401f
C11888 VDD.n4676 VSUBS 0.00283f
C11889 VDD.n4677 VSUBS 0.00307f
C11890 VDD.n4678 VSUBS 0.00134f
C11891 VDD.n4679 VSUBS 0.00201f
C11892 VDD.n4680 VSUBS 0.00378f
C11893 VDD.n4681 VSUBS 0.00134f
C11894 VDD.n4682 VSUBS 0.00741f
C11895 VDD.n4683 VSUBS 0.00194f
C11896 VDD.n4684 VSUBS 0.0198f
C11897 VDD.n4685 VSUBS 0.539f
C11898 VDD.n4686 VSUBS 0.509f
C11899 VDD.n4687 VSUBS 0.0155f
C11900 VDD.n4688 VSUBS 0.173f
C11901 VDD.n4689 VSUBS 0.183f
C11902 VDD.n4690 VSUBS 0.00661f
C11903 VDD.n4691 VSUBS 4.72e-19
C11904 VDD.n4692 VSUBS 0.00134f
C11905 VDD.n4693 VSUBS 0.00201f
C11906 VDD.n4694 VSUBS 0.00153f
C11907 VDD.n4695 VSUBS 0.00295f
C11908 VDD.n4696 VSUBS 0.00484f
C11909 VDD.n4697 VSUBS 0.00496f
C11910 VDD.n4698 VSUBS 0.00393f
C11911 VDD.n4699 VSUBS 0.00393f
C11912 VDD.n4700 VSUBS 0.00134f
C11913 VDD.n4701 VSUBS 0.00764f
C11914 VDD.n4702 VSUBS 0.00194f
C11915 VDD.n4703 VSUBS 0.0198f
C11916 VDD.n4704 VSUBS 0.539f
C11917 VDD.t15 VSUBS 0.366f
C11918 VDD.n4705 VSUBS 0.275f
C11919 VDD.n4706 VSUBS 0.0155f
C11920 VDD.n4707 VSUBS 0.173f
C11921 VDD.n4708 VSUBS 0.183f
C11922 VDD.n4709 VSUBS 0.00639f
C11923 VDD.n4710 VSUBS 4.72e-19
C11924 VDD.n4711 VSUBS 0.00134f
C11925 VDD.n4712 VSUBS 0.00201f
C11926 VDD.n4713 VSUBS 0.00106f
C11927 VDD.n4714 VSUBS 0.00271f
C11928 VDD.n4715 VSUBS 0.00496f
C11929 VDD.n4716 VSUBS 0.00354f
C11930 VDD.n4717 VSUBS 0.00409f
C11931 VDD.n4718 VSUBS 0.00248f
C11932 VDD.n4719 VSUBS 0.00409f
C11933 VDD.n4720 VSUBS 0.00134f
C11934 VDD.n4721 VSUBS 0.00593f
C11935 VDD.n4722 VSUBS 0.00194f
C11936 VDD.n4723 VSUBS 0.0198f
C11937 VDD.n4724 VSUBS 0.407f
C11938 VDD.n4725 VSUBS 0.509f
C11939 VDD.n4726 VSUBS 0.0155f
C11940 VDD.n4727 VSUBS 0.173f
C11941 VDD.n4728 VSUBS 0.183f
C11942 VDD.n4729 VSUBS 0.00616f
C11943 VDD.n4730 VSUBS 1.57e-19
C11944 VDD.n4731 VSUBS 0.00134f
C11945 VDD.n4732 VSUBS 0.00201f
C11946 VDD.n4733 VSUBS 0.0026f
C11947 VDD.n4734 VSUBS 0.00543f
C11948 VDD.n4735 VSUBS 0.00507f
C11949 VDD.n4736 VSUBS 0.00283f
C11950 VDD.n4737 VSUBS 8.26e-19
C11951 VDD.n4738 VSUBS 0.00409f
C11952 VDD.n4739 VSUBS 0.00134f
C11953 VDD.n4740 VSUBS 0.00593f
C11954 VDD.n4741 VSUBS 0.00194f
C11955 VDD.n4742 VSUBS 0.0198f
C11956 VDD.n4743 VSUBS 0.366f
C11957 VDD.n4744 VSUBS 0.183f
C11958 VDD.n4745 VSUBS 0.0155f
C11959 VDD.n4746 VSUBS 0.173f
C11960 VDD.n4747 VSUBS 0.499f
C11961 VDD.n4748 VSUBS 0.00616f
C11962 VDD.n4749 VSUBS 1.57e-19
C11963 VDD.n4750 VSUBS 0.00134f
C11964 VDD.n4751 VSUBS 0.00201f
C11965 VDD.n4752 VSUBS 0.00409f
C11966 VDD.n4753 VSUBS 0.00212f
C11967 VDD.n4754 VSUBS 0.00319f
C11968 VDD.n4755 VSUBS 0.0046f
C11969 VDD.n4756 VSUBS 0.00307f
C11970 VDD.n4757 VSUBS 0.00393f
C11971 VDD.n4758 VSUBS 0.00134f
C11972 VDD.n4759 VSUBS 0.00764f
C11973 VDD.n4760 VSUBS 0.00194f
C11974 VDD.t8 VSUBS 0.499f
C11975 VDD.n4761 VSUBS 0.0198f
C11976 VDD.n4762 VSUBS 0.0509f
C11977 VDD.n4763 VSUBS 0.183f
C11978 VDD.n4764 VSUBS 0.0155f
C11979 VDD.n4765 VSUBS 0.173f
C11980 VDD.n4766 VSUBS 0.509f
C11981 VDD.n4767 VSUBS 0.00639f
C11982 VDD.n4768 VSUBS 0.00157f
C11983 VDD.n4769 VSUBS 0.00342f
C11984 VDD.n4770 VSUBS 0.00417f
C11985 VDD.n4771 VSUBS 0.00496f
C11986 VDD.n4772 VSUBS 0.00413f
C11987 VDD.n4773 VSUBS 0.00307f
C11988 VDD.n4774 VSUBS 0.00378f
C11989 VDD.n4775 VSUBS 0.00118f
C11990 VDD.n4776 VSUBS 0.00741f
C11991 VDD.n4777 VSUBS 0.00194f
C11992 VDD.n4778 VSUBS 0.0198f
C11993 VDD.n4779 VSUBS 0.539f
C11994 VDD.n4780 VSUBS 0.183f
C11995 VDD.n4781 VSUBS 0.0155f
C11996 VDD.n4782 VSUBS 0.173f
C11997 VDD.n4783 VSUBS 0.509f
C11998 VDD.n4784 VSUBS 0.00661f
C11999 VDD.n4785 VSUBS 0.00126f
C12000 VDD.n4786 VSUBS 3.93e-19
C12001 VDD.n4787 VSUBS 0.00212f
C12002 VDD.n4788 VSUBS 0.00189f
C12003 VDD.n4789 VSUBS 0.00201f
C12004 VDD.n4790 VSUBS 8.26e-19
C12005 VDD.n4791 VSUBS 0.00134f
C12006 VDD.n4792 VSUBS 5.51e-19
C12007 VDD.n4793 VSUBS 0.00283f
C12008 VDD.n4794 VSUBS 0.00283f
C12009 VDD.n4795 VSUBS 0.00295f
C12010 VDD.n4796 VSUBS 0.00295f
C12011 VDD.n4797 VSUBS 0.0033f
C12012 VDD.n4798 VSUBS 0.00102f
C12013 VDD.n4799 VSUBS 0.00719f
C12014 VDD.n4800 VSUBS 0.00194f
C12015 VDD.n4801 VSUBS 0.0198f
C12016 VDD.n4802 VSUBS 0.539f
C12017 VDD.n4803 VSUBS 0.183f
C12018 VDD.n4804 VSUBS 0.0155f
C12019 VDD.n4805 VSUBS 0.132f
C12020 VDD.t2 VSUBS 0.0712f
C12021 VDD.n4806 VSUBS 0.478f
C12022 VDD.n4807 VSUBS 0.00684f
C12023 VDD.n4808 VSUBS 9.44e-19
C12024 VDD.n4809 VSUBS 5.51e-19
C12025 VDD.n4810 VSUBS 0.00283f
C12026 VDD.n4811 VSUBS 0.00142f
C12027 VDD.n4812 VSUBS 0.00201f
C12028 VDD.n4813 VSUBS 0.0013f
C12029 VDD.n4814 VSUBS 0.00134f
C12030 VDD.n4815 VSUBS 8.65e-19
C12031 VDD.n4816 VSUBS 0.00283f
C12032 VDD.n4817 VSUBS 0.00271f
C12033 VDD.n4818 VSUBS 0.00283f
C12034 VDD.n4819 VSUBS 0.00283f
C12035 VDD.n4820 VSUBS 0.0033f
C12036 VDD.n4821 VSUBS 8.65e-19
C12037 VDD.n4822 VSUBS 0.00134f
C12038 VDD.n4823 VSUBS 0.00696f
C12039 VDD.n4824 VSUBS 0.00194f
C12040 VDD.n4825 VSUBS 0.0198f
C12041 VDD.n4826 VSUBS 0.539f
C12042 VDD.n4827 VSUBS 0.183f
C12043 VDD.n4828 VSUBS 0.0155f
C12044 VDD.n4829 VSUBS 0.173f
C12045 VDD.n4830 VSUBS 0.0198f
C12046 VDD.n4831 VSUBS 0.539f
C12047 VDD.n4832 VSUBS 0.509f
C12048 VDD.n4833 VSUBS 0.00707f
C12049 VDD.n4834 VSUBS 6.29e-19
C12050 VDD.n4835 VSUBS 7.08e-19
C12051 VDD.n4836 VSUBS 0.00319f
C12052 VDD.n4837 VSUBS 9.44e-19
C12053 VDD.n4838 VSUBS 0.00201f
C12054 VDD.n4839 VSUBS 0.00401f
C12055 VDD.n4840 VSUBS 0.00378f
C12056 VDD.n4841 VSUBS 0.00307f
C12057 VDD.n4842 VSUBS 0.00401f
C12058 VDD.n4843 VSUBS 0.0033f
C12059 VDD.n4844 VSUBS 0.00118f
C12060 VDD.n4845 VSUBS 8.65e-19
C12061 VDD.n4846 VSUBS 0.00319f
C12062 VDD.n4847 VSUBS 0.00201f
C12063 VDD.n4848 VSUBS 0.00673f
C12064 VDD.n4849 VSUBS 0.00194f
C12065 VDD.n4850 VSUBS 0.183f
C12066 VDD.n4851 VSUBS 0.0155f
C12067 VDD.n4852 VSUBS 0.173f
C12068 VDD.t187 VSUBS 0.397f
C12069 VDD.n4853 VSUBS 0.254f
C12070 VDD.n4854 VSUBS 0.0073f
C12071 VDD.n4855 VSUBS 0.00134f
C12072 VDD.n4856 VSUBS 0.00299f
C12073 VDD.n4857 VSUBS 0.00134f
C12074 VDD.n4858 VSUBS 0.00201f
C12075 VDD.n4859 VSUBS 0.00153f
C12076 VDD.n4860 VSUBS 0.00283f
C12077 VDD.n4861 VSUBS 0.00496f
C12078 VDD.n4862 VSUBS 0.00496f
C12079 VDD.n4863 VSUBS 0.00315f
C12080 VDD.n4864 VSUBS 0.00134f
C12081 VDD.n4865 VSUBS 0.0065f
C12082 VDD.n4866 VSUBS 0.00194f
C12083 VDD.n4867 VSUBS 0.0198f
C12084 VDD.n4868 VSUBS 0.397f
C12085 VDD.n4869 VSUBS 0.183f
C12086 VDD.n4870 VSUBS 0.0155f
C12087 VDD.n4871 VSUBS 0.173f
C12088 VDD.n4872 VSUBS 0.509f
C12089 VDD.n4873 VSUBS 0.00753f
C12090 VDD.n4874 VSUBS 0.00205f
C12091 VDD.n4875 VSUBS 0.00315f
C12092 VDD.n4876 VSUBS 0.00134f
C12093 VDD.n4877 VSUBS 0.00201f
C12094 VDD.n4878 VSUBS 0.00106f
C12095 VDD.n4879 VSUBS 0.0026f
C12096 VDD.n4880 VSUBS 0.00496f
C12097 VDD.n4881 VSUBS 0.00366f
C12098 VDD.n4882 VSUBS 0.00248f
C12099 VDD.n4883 VSUBS 0.00299f
C12100 VDD.n4884 VSUBS 0.00134f
C12101 VDD.n4885 VSUBS 0.00627f
C12102 VDD.n4886 VSUBS 0.00194f
C12103 VDD.n4887 VSUBS 0.0198f
C12104 VDD.n4888 VSUBS 0.539f
C12105 VDD.n4889 VSUBS 0.183f
C12106 VDD.n4890 VSUBS 0.0155f
C12107 VDD.n4891 VSUBS 0.173f
C12108 VDD.n4892 VSUBS 0.0155f
C12109 VDD.n4893 VSUBS 0.692f
C12110 VDD.n4894 VSUBS 0.0198f
C12111 VDD.n4895 VSUBS 0.214f
C12112 VDD.t83 VSUBS 0.356f
C12113 VDD.n4896 VSUBS 0.478f
C12114 VDD.n4897 VSUBS 0.00776f
C12115 VDD.n4898 VSUBS 0.00236f
C12116 VDD.n4899 VSUBS 0.00299f
C12117 VDD.n4900 VSUBS 0.00134f
C12118 VDD.n4901 VSUBS 0.00189f
C12119 VDD.n4902 VSUBS 2.36e-19
C12120 VDD.n4903 VSUBS 0.00248f
C12121 VDD.n4904 VSUBS 0.00531f
C12122 VDD.n4905 VSUBS 0.00507f
C12123 VDD.n4906 VSUBS 0.00295f
C12124 VDD.n4907 VSUBS 0.0138f
C12125 VDD.n4908 VSUBS 0.00551f
C12126 VDD.n4909 VSUBS 0.0138f
C12127 VDD.n4910 VSUBS 0.00543f
C12128 VDD.n4911 VSUBS 0.00535f
C12129 VDD.n4912 VSUBS 0.00295f
C12130 VDD.n4913 VSUBS 0.00507f
C12131 VDD.n4914 VSUBS 0.0046f
C12132 VDD.n4915 VSUBS 0.00307f
C12133 VDD.n4916 VSUBS 0.00134f
C12134 VDD.n4917 VSUBS 0.00283f
C12135 VDD.n4918 VSUBS 0.00153f
C12136 VDD.n4919 VSUBS 0.00201f
C12137 VDD.n4920 VSUBS 0.00134f
C12138 VDD.n4921 VSUBS 0.00201f
C12139 VDD.n4922 VSUBS 0.00275f
C12140 VDD.n4923 VSUBS 0.00134f
C12141 VDD.n4924 VSUBS 0.00627f
C12142 VDD.n4925 VSUBS 0.00194f
C12143 VDD.n4926 VSUBS 0.0198f
C12144 VDD.n4927 VSUBS 0.692f
C12145 VDD.n4928 VSUBS 0.0155f
C12146 VDD.n4929 VSUBS 0.692f
C12147 VDD.n4930 VSUBS 0.0198f
C12148 VDD.n4931 VSUBS 0.539f
C12149 VDD.n4932 VSUBS 0.499f
C12150 VDD.t98 VSUBS 0.0203f
C12151 VDD.n4933 VSUBS 0.0155f
C12152 VDD.n4934 VSUBS 0.163f
C12153 VDD.n4935 VSUBS 0.183f
C12154 VDD.n4936 VSUBS 0.00776f
C12155 VDD.n4937 VSUBS 0.00126f
C12156 VDD.n4938 VSUBS 0.00295f
C12157 VDD.n4939 VSUBS 0.00401f
C12158 VDD.n4940 VSUBS 0.00307f
C12159 VDD.n4941 VSUBS 0.00126f
C12160 VDD.n4942 VSUBS 0.00283f
C12161 VDD.n4943 VSUBS 0.00224f
C12162 VDD.n4944 VSUBS 0.00189f
C12163 VDD.n4945 VSUBS 0.00201f
C12164 VDD.n4946 VSUBS 8.26e-19
C12165 VDD.n4947 VSUBS 0.00134f
C12166 VDD.n4948 VSUBS 0.0065f
C12167 VDD.n4949 VSUBS 0.00194f
C12168 VDD.n4950 VSUBS 0.0198f
C12169 VDD.n4951 VSUBS 0.539f
C12170 VDD.n4952 VSUBS 0.509f
C12171 VDD.n4953 VSUBS 0.0155f
C12172 VDD.n4954 VSUBS 0.173f
C12173 VDD.n4955 VSUBS 0.183f
C12174 VDD.n4956 VSUBS 0.00753f
C12175 VDD.n4957 VSUBS 5.51e-19
C12176 VDD.n4958 VSUBS 0.00275f
C12177 VDD.n4959 VSUBS 0.0011f
C12178 VDD.n4960 VSUBS 0.00102f
C12179 VDD.n4961 VSUBS 0.00271f
C12180 VDD.n4962 VSUBS 0.00295f
C12181 VDD.n4963 VSUBS 0.00295f
C12182 VDD.n4964 VSUBS 9.44e-19
C12183 VDD.n4965 VSUBS 0.00283f
C12184 VDD.n4966 VSUBS 0.00295f
C12185 VDD.n4967 VSUBS 0.00142f
C12186 VDD.n4968 VSUBS 0.00201f
C12187 VDD.n4969 VSUBS 0.0013f
C12188 VDD.n4970 VSUBS 0.00134f
C12189 VDD.n4971 VSUBS 0.00673f
C12190 VDD.n4972 VSUBS 0.00194f
C12191 VDD.n4973 VSUBS 0.0198f
C12192 VDD.n4974 VSUBS 0.539f
C12193 VDD.t76 VSUBS 0.448f
C12194 VDD.n4975 VSUBS 0.234f
C12195 VDD.n4976 VSUBS 0.0155f
C12196 VDD.n4977 VSUBS 0.173f
C12197 VDD.n4978 VSUBS 0.183f
C12198 VDD.n4979 VSUBS 0.0073f
C12199 VDD.n4980 VSUBS 8.65e-19
C12200 VDD.n4981 VSUBS 0.00275f
C12201 VDD.n4982 VSUBS 0.00126f
C12202 VDD.n4983 VSUBS 8.65e-19
C12203 VDD.n4984 VSUBS 0.0026f
C12204 VDD.n4985 VSUBS 0.00283f
C12205 VDD.n4986 VSUBS 0.00283f
C12206 VDD.n4987 VSUBS 0.00126f
C12207 VDD.n4988 VSUBS 6.29e-19
C12208 VDD.n4989 VSUBS 0.00283f
C12209 VDD.n4990 VSUBS 0.0033f
C12210 VDD.n4991 VSUBS 9.44e-19
C12211 VDD.n4992 VSUBS 0.00189f
C12212 VDD.n4993 VSUBS 0.00322f
C12213 VDD.n4994 VSUBS 0.00134f
C12214 VDD.n4995 VSUBS 0.00696f
C12215 VDD.n4996 VSUBS 0.00194f
C12216 VDD.n4997 VSUBS 0.0198f
C12217 VDD.n4998 VSUBS 0.366f
C12218 VDD.n4999 VSUBS 0.509f
C12219 VDD.n5000 VSUBS 0.0155f
C12220 VDD.n5001 VSUBS 0.173f
C12221 VDD.n5002 VSUBS 0.183f
C12222 VDD.n5003 VSUBS 0.00707f
C12223 VDD.n5004 VSUBS 7.87e-19
C12224 VDD.n5005 VSUBS 0.00126f
C12225 VDD.n5006 VSUBS 0.00189f
C12226 VDD.n5007 VSUBS 0.00201f
C12227 VDD.n5008 VSUBS 0.00295f
C12228 VDD.n5009 VSUBS 0.00401f
C12229 VDD.n5010 VSUBS 0.00283f
C12230 VDD.n5011 VSUBS 0.0033f
C12231 VDD.n5012 VSUBS 0.00201f
C12232 VDD.n5013 VSUBS 0.00134f
C12233 VDD.n5014 VSUBS 0.00362f
C12234 VDD.n5015 VSUBS 0.00134f
C12235 VDD.n5016 VSUBS 0.00719f
C12236 VDD.n5017 VSUBS 0.00194f
C12237 VDD.n5018 VSUBS 0.0198f
C12238 VDD.n5019 VSUBS 0.539f
C12239 VDD.n5020 VSUBS 0.458f
C12240 VDD.n5021 VSUBS 0.0155f
C12241 VDD.n5022 VSUBS 0.173f
C12242 VDD.n5023 VSUBS 0.183f
C12243 VDD.n5024 VSUBS 0.00684f
C12244 VDD.n5025 VSUBS 7.87e-19
C12245 VDD.n5026 VSUBS 0.00134f
C12246 VDD.n5027 VSUBS 0.00201f
C12247 VDD.n5028 VSUBS 0.00153f
C12248 VDD.n5029 VSUBS 0.00271f
C12249 VDD.n5030 VSUBS 0.00507f
C12250 VDD.n5031 VSUBS 0.00496f
C12251 VDD.n5032 VSUBS 0.00378f
C12252 VDD.n5033 VSUBS 0.00378f
C12253 VDD.n5034 VSUBS 0.00134f
C12254 VDD.n5035 VSUBS 0.00741f
C12255 VDD.n5036 VSUBS 0.00194f
C12256 VDD.t117 VSUBS 0.407f
C12257 VDD.n5037 VSUBS 0.0198f
C12258 VDD.n5038 VSUBS 0.183f
C12259 VDD.n5039 VSUBS 0.509f
C12260 VDD.n5040 VSUBS 0.0155f
C12261 VDD.n5041 VSUBS 0.173f
C12262 VDD.n5042 VSUBS 0.183f
C12263 VDD.n5043 VSUBS 0.00661f
C12264 VDD.n5044 VSUBS 7.87e-19
C12265 VDD.n5045 VSUBS 0.00134f
C12266 VDD.n5046 VSUBS 0.00201f
C12267 VDD.n5047 VSUBS 0.00106f
C12268 VDD.n5048 VSUBS 0.00248f
C12269 VDD.n5049 VSUBS 0.00496f
C12270 VDD.n5050 VSUBS 0.00378f
C12271 VDD.n5051 VSUBS 0.00248f
C12272 VDD.n5052 VSUBS 0.00393f
C12273 VDD.n5053 VSUBS 0.00393f
C12274 VDD.n5054 VSUBS 0.00134f
C12275 VDD.n5055 VSUBS 0.00764f
C12276 VDD.n5056 VSUBS 0.00194f
C12277 VDD.n5057 VSUBS 0.0198f
C12278 VDD.n5058 VSUBS 0.539f
C12279 VDD.n5059 VSUBS 0.509f
C12280 VDD.n5060 VSUBS 0.0155f
C12281 VDD.n5061 VSUBS 0.173f
C12282 VDD.n5062 VSUBS 0.183f
C12283 VDD.n5063 VSUBS 0.00639f
C12284 VDD.n5064 VSUBS 4.72e-19
C12285 VDD.n5065 VSUBS 0.00134f
C12286 VDD.n5066 VSUBS 0.00177f
C12287 VDD.n5067 VSUBS 3.54e-19
C12288 VDD.n5068 VSUBS 0.00248f
C12289 VDD.n5069 VSUBS 0.00519f
C12290 VDD.n5070 VSUBS 0.00401f
C12291 VDD.n5071 VSUBS 0.00409f
C12292 VDD.n5072 VSUBS 0.00212f
C12293 VDD.n5073 VSUBS 0.00189f
C12294 VDD.n5074 VSUBS 0.00409f
C12295 VDD.n5075 VSUBS 0.00134f
C12296 VDD.n5076 VSUBS 0.00593f
C12297 VDD.n5077 VSUBS 0.00194f
C12298 VDD.n5078 VSUBS 0.539f
C12299 VDD.n5079 VSUBS 0.509f
C12300 VDD.n5080 VSUBS 0.0155f
C12301 VDD.n5081 VSUBS 0.173f
C12302 VDD.t120 VSUBS 0.183f
C12303 VDD.n5082 VSUBS 0.00616f
C12304 VDD.n5083 VSUBS 1.57e-19
C12305 VDD.n5084 VSUBS 0.00134f
C12306 VDD.n5085 VSUBS 9.44e-19
C12307 VDD.n5086 VSUBS 0.00212f
C12308 VDD.n5087 VSUBS 0.00496f
C12309 VDD.n5088 VSUBS 0.0046f
C12310 VDD.n5089 VSUBS 0.00307f
C12311 VDD.n5090 VSUBS 0.00401f
C12312 VDD.n5091 VSUBS 0.00593f
C12313 VDD.n5092 VSUBS 0.00194f
C12314 VDD.n5093 VSUBS 0.366f
C12315 VDD.n5094 VSUBS 0.183f
C12316 VDD.n5095 VSUBS 0.173f
C12317 VDD.n5096 VSUBS 0.509f
C12318 VDD.n5097 VSUBS 0.00616f
C12319 VDD.n5098 VSUBS 0.00126f
C12320 VDD.n5099 VSUBS 1.57e-19
C12321 VDD.n5100 VSUBS 0.00126f
C12322 VDD.n5101 VSUBS 0.00165f
C12323 VDD.n5102 VSUBS 0.00201f
C12324 VDD.n5103 VSUBS 0.00134f
C12325 VDD.n5104 VSUBS 0.00201f
C12326 VDD.n5105 VSUBS 0.00299f
C12327 VDD.n5106 VSUBS 0.00295f
C12328 VDD.n5107 VSUBS 0.00389f
C12329 VDD.n5108 VSUBS 0.00307f
C12330 VDD.n5109 VSUBS 0.00385f
C12331 VDD.n5110 VSUBS 0.00764f
C12332 VDD.n5111 VSUBS 0.00194f
C12333 VDD.n5112 VSUBS 0.539f
C12334 VDD.n5113 VSUBS 0.183f
C12335 VDD.n5114 VSUBS 0.173f
C12336 VDD.t24 VSUBS 0.478f
C12337 VDD.n5115 VSUBS 0.214f
C12338 VDD.n5116 VSUBS 0.00639f
C12339 VDD.n5117 VSUBS 0.00118f
C12340 VDD.n5118 VSUBS 3.15e-19
C12341 VDD.n5119 VSUBS 0.0011f
C12342 VDD.n5120 VSUBS 0.00236f
C12343 VDD.n5121 VSUBS 0.00189f
C12344 VDD.n5122 VSUBS 0.00201f
C12345 VDD.n5123 VSUBS 8.26e-19
C12346 VDD.n5124 VSUBS 0.00134f
C12347 VDD.n5125 VSUBS 5.51e-19
C12348 VDD.n5126 VSUBS 0.00283f
C12349 VDD.n5127 VSUBS 0.0026f
C12350 VDD.n5128 VSUBS 0.00295f
C12351 VDD.n5129 VSUBS 0.00295f
C12352 VDD.n5130 VSUBS 0.00354f
C12353 VDD.n5131 VSUBS 0.00741f
C12354 VDD.n5132 VSUBS 0.00194f
C12355 VDD.n5133 VSUBS 0.356f
C12356 VDD.n5134 VSUBS 0.183f
C12357 VDD.n5135 VSUBS 0.173f
C12358 VDD.n5136 VSUBS 0.509f
C12359 VDD.n5137 VSUBS 0.00661f
C12360 VDD.n5138 VSUBS 8.65e-19
C12361 VDD.n5139 VSUBS 4.72e-19
C12362 VDD.n5140 VSUBS 9.44e-19
C12363 VDD.n5141 VSUBS 0.00307f
C12364 VDD.n5142 VSUBS 0.00142f
C12365 VDD.n5143 VSUBS 0.00201f
C12366 VDD.n5144 VSUBS 0.00134f
C12367 VDD.n5145 VSUBS 0.0037f
C12368 VDD.n5146 VSUBS 0.00378f
C12369 VDD.n5147 VSUBS 0.00283f
C12370 VDD.n5148 VSUBS 0.00283f
C12371 VDD.n5149 VSUBS 0.00354f
C12372 VDD.n5150 VSUBS 6.29e-19
C12373 VDD.n5151 VSUBS 7.87e-19
C12374 VDD.n5152 VSUBS 0.00342f
C12375 VDD.n5153 VSUBS 0.00719f
C12376 VDD.n5154 VSUBS 0.00194f
C12377 VDD.n5155 VSUBS 0.0378f
C12378 VDD.n5156 VSUBS 0.539f
C12379 VDD.n5157 VSUBS 0.183f
C12380 VDD.n5158 VSUBS 0.173f
C12381 VDD.n5159 VSUBS 0.0595f
C12382 VDD.n5195 VSUBS 2.65f
C12383 VDD.n5196 VSUBS 0.801f
C12384 VDD.n5197 VSUBS 0.926f
C12385 VDD.n5198 VSUBS 1.38f
C12386 VDD.n5199 VSUBS 1.38f
C12387 VDD.n5200 VSUBS 0.895f
C12388 VDD.n5261 VSUBS 0.692f
C12389 VDD.n5262 VSUBS 0.926f
C12390 VDD.n5263 VSUBS 0.509f
C12391 VDD.n5264 VSUBS 0.0112f
C12392 VDD.n5265 VSUBS 0.00173f
C12393 VDD.n5266 VSUBS 0.00271f
C12394 VDD.n5267 VSUBS 0.00464f
C12395 VDD.n5268 VSUBS 0.00134f
C12396 VDD.n5269 VSUBS 0.00201f
C12397 VDD.n5270 VSUBS 0.00201f
C12398 VDD.n5271 VSUBS 0.0155f
C12399 VDD.n5272 VSUBS 0.0448f
C12400 VDD.n5273 VSUBS 0.0198f
C12401 VDD.n5274 VSUBS 0.0448f
C12402 VDD.n5275 VSUBS 0.0181f
C12403 VDD.n5276 VSUBS 0.0448f
C12404 VDD.n5277 VSUBS 0.0198f
C12405 VDD.n5278 VSUBS 0.0494f
C12406 VDD.n5279 VSUBS 0.0198f
C12407 VDD.n5280 VSUBS 0.0744f
C12408 VDD.n5281 VSUBS 0.0198f
C12409 VDD.n5282 VSUBS 0.0448f
C12410 VDD.n5283 VSUBS 0.0155f
C12411 VDD.n5284 VSUBS 0.0448f
C12412 VDD.n5285 VSUBS 0.0198f
C12413 VDD.n5286 VSUBS 0.0448f
C12414 VDD.n5287 VSUBS 0.0155f
C12415 VDD.n5288 VSUBS 0.0448f
C12416 VDD.n5289 VSUBS 0.0198f
C12417 VDD.n5290 VSUBS 0.0448f
C12418 VDD.n5291 VSUBS 0.0155f
C12419 VDD.n5292 VSUBS 0.0448f
C12420 VDD.n5293 VSUBS 0.0198f
C12421 VDD.n5294 VSUBS 0.0448f
C12422 VDD.n5295 VSUBS 0.0155f
C12423 VDD.n5296 VSUBS 0.0448f
C12424 VDD.n5297 VSUBS 0.0198f
C12425 VDD.n5298 VSUBS 0.0448f
C12426 VDD.n5299 VSUBS 0.0155f
C12427 VDD.n5300 VSUBS 0.0448f
C12428 VDD.n5301 VSUBS 0.0198f
C12429 VDD.n5302 VSUBS 0.0448f
C12430 VDD.n5303 VSUBS 0.0155f
C12431 VDD.n5304 VSUBS 0.0448f
C12432 VDD.n5305 VSUBS 0.0198f
C12433 VDD.n5306 VSUBS 0.0448f
C12434 VDD.n5307 VSUBS 0.0155f
C12435 VDD.n5308 VSUBS 0.0448f
C12436 VDD.n5309 VSUBS 0.0198f
C12437 VDD.n5310 VSUBS 0.0448f
C12438 VDD.n5311 VSUBS 0.0155f
C12439 VDD.n5312 VSUBS 0.0448f
C12440 VDD.n5313 VSUBS 0.0198f
C12441 VDD.n5314 VSUBS 0.0448f
C12442 VDD.n5315 VSUBS 0.0155f
C12443 VDD.n5316 VSUBS 0.0448f
C12444 VDD.n5317 VSUBS 0.0198f
C12445 VDD.n5318 VSUBS 0.0448f
C12446 VDD.n5319 VSUBS 0.0155f
C12447 VDD.n5320 VSUBS 0.0448f
C12448 VDD.n5321 VSUBS 0.0198f
C12449 VDD.n5322 VSUBS 0.0448f
C12450 VDD.n5323 VSUBS 0.0155f
C12451 VDD.n5324 VSUBS 0.0448f
C12452 VDD.n5325 VSUBS 0.0198f
C12453 VDD.n5326 VSUBS 0.0448f
C12454 VDD.n5327 VSUBS 0.0155f
C12455 VDD.n5328 VSUBS 0.0448f
C12456 VDD.n5329 VSUBS 0.0198f
C12457 VDD.n5330 VSUBS 0.0448f
C12458 VDD.n5331 VSUBS 0.0155f
C12459 VDD.n5332 VSUBS 0.0448f
C12460 VDD.n5333 VSUBS 0.0198f
C12461 VDD.n5334 VSUBS 0.0448f
C12462 VDD.n5335 VSUBS 0.0155f
C12463 VDD.n5336 VSUBS 0.0448f
C12464 VDD.n5337 VSUBS 0.0198f
C12465 VDD.n5338 VSUBS 0.0448f
C12466 VDD.n5339 VSUBS 0.0155f
C12467 VDD.n5340 VSUBS 0.0448f
C12468 VDD.n5341 VSUBS 0.0198f
C12469 VDD.n5342 VSUBS 0.0448f
C12470 VDD.n5343 VSUBS 0.0155f
C12471 VDD.n5344 VSUBS 0.0448f
C12472 VDD.n5345 VSUBS 0.0198f
C12473 VDD.n5346 VSUBS 0.0448f
C12474 VDD.n5347 VSUBS 0.0181f
C12475 VDD.n5348 VSUBS 0.0448f
C12476 VDD.n5349 VSUBS 0.0198f
C12477 VDD.n5350 VSUBS 0.0639f
C12478 VDD.n5351 VSUBS 0.0198f
C12479 VDD.n5352 VSUBS 0.0599f
C12480 VDD.n5353 VSUBS 0.0495f
C12481 VDD.n5354 VSUBS 0.019f
C12482 VDD.n5355 VSUBS 0.00283f
C12483 VDD.n5356 VSUBS 0.00307f
C12484 VDD.n5357 VSUBS 0.00661f
C12485 VDD.n5358 VSUBS 0.00763f
C12486 VDD.n5359 VSUBS 0.00397f
C12487 VDD.n5360 VSUBS 0.0145f
C12488 VDD.t380 VSUBS 0.0114f
C12489 VDD.t63 VSUBS 0.0114f
C12490 VDD.n5361 VSUBS 0.0267f
C12491 VDD.n5362 VSUBS 0.0114f
C12492 VDD.n5363 VSUBS 0.0229f
C12493 VDD.n5364 VSUBS 0.0142f
C12494 VDD.n5365 VSUBS 0.00763f
C12495 VDD.n5366 VSUBS 0.00397f
C12496 VDD.n5367 VSUBS 0.0145f
C12497 VDD.t411 VSUBS 0.0114f
C12498 VDD.t389 VSUBS 0.0114f
C12499 VDD.n5368 VSUBS 0.0267f
C12500 VDD.n5369 VSUBS 0.0114f
C12501 VDD.n5370 VSUBS 0.0229f
C12502 VDD.n5371 VSUBS 0.0142f
C12503 VDD.n5372 VSUBS 0.00763f
C12504 VDD.n5373 VSUBS 0.00397f
C12505 VDD.n5374 VSUBS 0.0145f
C12506 VDD.t443 VSUBS 0.0114f
C12507 VDD.t99 VSUBS 0.0114f
C12508 VDD.n5375 VSUBS 0.0267f
C12509 VDD.n5376 VSUBS 0.0114f
C12510 VDD.n5377 VSUBS 0.0229f
C12511 VDD.n5378 VSUBS 0.0142f
C12512 VDD.n5379 VSUBS 0.00763f
C12513 VDD.n5380 VSUBS 0.00397f
C12514 VDD.n5381 VSUBS 0.0145f
C12515 VDD.t378 VSUBS 0.0114f
C12516 VDD.t408 VSUBS 0.0114f
C12517 VDD.n5382 VSUBS 0.0267f
C12518 VDD.n5383 VSUBS 0.0114f
C12519 VDD.n5384 VSUBS 0.0229f
C12520 VDD.n5385 VSUBS 0.0142f
C12521 VDD.n5386 VSUBS 0.00763f
C12522 VDD.n5387 VSUBS 0.00397f
C12523 VDD.n5388 VSUBS 0.0145f
C12524 VDD.t52 VSUBS 0.0114f
C12525 VDD.t68 VSUBS 0.0114f
C12526 VDD.n5389 VSUBS 0.0267f
C12527 VDD.n5390 VSUBS 0.0114f
C12528 VDD.n5391 VSUBS 0.0229f
C12529 VDD.n5392 VSUBS 0.0142f
C12530 VDD.n5393 VSUBS 0.00763f
C12531 VDD.n5394 VSUBS 0.00397f
C12532 VDD.n5395 VSUBS 0.0145f
C12533 VDD.t394 VSUBS 0.0114f
C12534 VDD.t405 VSUBS 0.0114f
C12535 VDD.n5396 VSUBS 0.0267f
C12536 VDD.n5397 VSUBS 0.0114f
C12537 VDD.n5398 VSUBS 0.0229f
C12538 VDD.n5399 VSUBS 0.0142f
C12539 VDD.n5400 VSUBS 0.00763f
C12540 VDD.n5401 VSUBS 0.00397f
C12541 VDD.n5402 VSUBS 0.0145f
C12542 VDD.t465 VSUBS 0.0114f
C12543 VDD.t22 VSUBS 0.0114f
C12544 VDD.n5403 VSUBS 0.0267f
C12545 VDD.n5404 VSUBS 0.0114f
C12546 VDD.n5405 VSUBS 0.0229f
C12547 VDD.n5406 VSUBS 0.0142f
C12548 VDD.n5407 VSUBS 0.00763f
C12549 VDD.n5408 VSUBS 0.00397f
C12550 VDD.n5409 VSUBS 0.0145f
C12551 VDD.t71 VSUBS 0.0114f
C12552 VDD.t428 VSUBS 0.0114f
C12553 VDD.n5410 VSUBS 0.0267f
C12554 VDD.n5411 VSUBS 0.0114f
C12555 VDD.n5412 VSUBS 0.0229f
C12556 VDD.n5413 VSUBS 0.0142f
C12557 VDD.n5414 VSUBS 0.00763f
C12558 VDD.n5415 VSUBS 0.00397f
C12559 VDD.n5416 VSUBS 0.0145f
C12560 VDD.t79 VSUBS 0.0114f
C12561 VDD.t153 VSUBS 0.0114f
C12562 VDD.n5417 VSUBS 0.0267f
C12563 VDD.n5418 VSUBS 0.0114f
C12564 VDD.n5419 VSUBS 0.0229f
C12565 VDD.n5420 VSUBS 0.0142f
C12566 VDD.n5421 VSUBS 0.00763f
C12567 VDD.n5422 VSUBS 0.00397f
C12568 VDD.n5423 VSUBS 0.0145f
C12569 VDD.t14 VSUBS 0.0114f
C12570 VDD.t466 VSUBS 0.0114f
C12571 VDD.n5424 VSUBS 0.0267f
C12572 VDD.n5425 VSUBS 0.0114f
C12573 VDD.n5426 VSUBS 0.0229f
C12574 VDD.n5427 VSUBS 0.0142f
C12575 VDD.n5428 VSUBS 0.00763f
C12576 VDD.n5429 VSUBS 0.00397f
C12577 VDD.n5430 VSUBS 0.0145f
C12578 VDD.t142 VSUBS 0.0114f
C12579 VDD.t167 VSUBS 0.0114f
C12580 VDD.n5431 VSUBS 0.0267f
C12581 VDD.n5432 VSUBS 0.0114f
C12582 VDD.n5433 VSUBS 0.0229f
C12583 VDD.n5434 VSUBS 0.0142f
C12584 VDD.n5435 VSUBS 0.00763f
C12585 VDD.n5436 VSUBS 0.00397f
C12586 VDD.n5437 VSUBS 0.0145f
C12587 VDD.t461 VSUBS 0.0114f
C12588 VDD.t423 VSUBS 0.0114f
C12589 VDD.n5438 VSUBS 0.0267f
C12590 VDD.n5439 VSUBS 0.0114f
C12591 VDD.n5440 VSUBS 0.0229f
C12592 VDD.n5441 VSUBS 0.0142f
C12593 VDD.n5442 VSUBS 0.00763f
C12594 VDD.n5443 VSUBS 0.00397f
C12595 VDD.n5444 VSUBS 0.0145f
C12596 VDD.t419 VSUBS 0.0114f
C12597 VDD.t141 VSUBS 0.0114f
C12598 VDD.n5445 VSUBS 0.0267f
C12599 VDD.n5446 VSUBS 0.0114f
C12600 VDD.n5447 VSUBS 0.0229f
C12601 VDD.n5448 VSUBS 0.0142f
C12602 VDD.n5449 VSUBS 0.00763f
C12603 VDD.n5450 VSUBS 0.00397f
C12604 VDD.n5451 VSUBS 0.0145f
C12605 VDD.t444 VSUBS 0.0114f
C12606 VDD.t127 VSUBS 0.0114f
C12607 VDD.n5452 VSUBS 0.0267f
C12608 VDD.n5453 VSUBS 0.0114f
C12609 VDD.n5454 VSUBS 0.0229f
C12610 VDD.n5455 VSUBS 0.0142f
C12611 VDD.n5456 VSUBS 0.00763f
C12612 VDD.n5457 VSUBS 0.00397f
C12613 VDD.n5458 VSUBS 0.0145f
C12614 VDD.t435 VSUBS 0.0114f
C12615 VDD.t152 VSUBS 0.0114f
C12616 VDD.n5459 VSUBS 0.0267f
C12617 VDD.n5460 VSUBS 0.0114f
C12618 VDD.n5461 VSUBS 0.0229f
C12619 VDD.n5462 VSUBS 0.0142f
C12620 VDD.n5463 VSUBS 0.00763f
C12621 VDD.n5464 VSUBS 0.00397f
C12622 VDD.n5465 VSUBS 0.0145f
C12623 VDD.t81 VSUBS 0.0114f
C12624 VDD.t391 VSUBS 0.0114f
C12625 VDD.n5466 VSUBS 0.0267f
C12626 VDD.n5467 VSUBS 0.0114f
C12627 VDD.n5468 VSUBS 0.0229f
C12628 VDD.n5469 VSUBS 0.0142f
C12629 VDD.n5470 VSUBS 0.00763f
C12630 VDD.n5471 VSUBS 0.00397f
C12631 VDD.n5472 VSUBS 0.0145f
C12632 VDD.t18 VSUBS 0.0114f
C12633 VDD.t397 VSUBS 0.0114f
C12634 VDD.n5473 VSUBS 0.0267f
C12635 VDD.n5474 VSUBS 0.0114f
C12636 VDD.n5475 VSUBS 0.0229f
C12637 VDD.n5476 VSUBS 0.0142f
C12638 VDD.n5477 VSUBS 0.00763f
C12639 VDD.n5478 VSUBS 0.00397f
C12640 VDD.n5479 VSUBS 0.0145f
C12641 VDD.t436 VSUBS 0.0114f
C12642 VDD.t100 VSUBS 0.0114f
C12643 VDD.n5480 VSUBS 0.0267f
C12644 VDD.n5481 VSUBS 0.0114f
C12645 VDD.n5482 VSUBS 0.0229f
C12646 VDD.n5483 VSUBS 0.0142f
C12647 VDD.n5484 VSUBS 0.00763f
C12648 VDD.n5485 VSUBS 0.00397f
C12649 VDD.n5486 VSUBS 0.0145f
C12650 VDD.t165 VSUBS 0.0114f
C12651 VDD.t458 VSUBS 0.0114f
C12652 VDD.n5487 VSUBS 0.0267f
C12653 VDD.n5488 VSUBS 0.0114f
C12654 VDD.n5489 VSUBS 0.0229f
C12655 VDD.n5490 VSUBS 0.0142f
C12656 VDD.n5491 VSUBS 0.00763f
C12657 VDD.n5492 VSUBS 0.00397f
C12658 VDD.n5493 VSUBS 0.0202f
C12659 VDD.t456 VSUBS 0.0114f
C12660 VDD.t414 VSUBS 0.0114f
C12661 VDD.n5494 VSUBS 0.0267f
C12662 VDD.n5495 VSUBS 0.0114f
C12663 VDD.n5496 VSUBS 0.0229f
C12664 VDD.n5497 VSUBS 0.0142f
C12665 VDD.n5498 VSUBS 0.215f
C12666 VDD.n5499 VSUBS 0.0867f
C12667 VDD.n5500 VSUBS 0.0867f
C12668 VDD.n5501 VSUBS 0.0867f
C12669 VDD.n5502 VSUBS 0.0867f
C12670 VDD.n5503 VSUBS 0.0867f
C12671 VDD.n5504 VSUBS 0.0867f
C12672 VDD.n5505 VSUBS 0.0867f
C12673 VDD.n5506 VSUBS 0.0867f
C12674 VDD.n5507 VSUBS 0.0867f
C12675 VDD.n5508 VSUBS 0.0867f
C12676 VDD.n5509 VSUBS 0.0867f
C12677 VDD.n5510 VSUBS 0.0867f
C12678 VDD.n5511 VSUBS 0.0867f
C12679 VDD.n5512 VSUBS 0.0867f
C12680 VDD.n5513 VSUBS 0.0867f
C12681 VDD.n5514 VSUBS 0.0867f
C12682 VDD.n5515 VSUBS 0.0867f
C12683 VDD.n5516 VSUBS 0.0867f
C12684 VDD.n5517 VSUBS 0.0867f
C12685 VDD.n5518 VSUBS 0.0867f
C12686 VDD.n5519 VSUBS 0.0867f
C12687 VDD.n5520 VSUBS 0.0867f
C12688 VDD.n5521 VSUBS 0.0867f
C12689 VDD.n5522 VSUBS 0.0867f
C12690 VDD.n5523 VSUBS 0.0867f
C12691 VDD.n5524 VSUBS 0.0867f
C12692 VDD.n5525 VSUBS 0.0867f
C12693 VDD.n5526 VSUBS 0.0867f
C12694 VDD.n5527 VSUBS 0.0867f
C12695 VDD.n5528 VSUBS 0.0867f
C12696 VDD.n5529 VSUBS 0.0867f
C12697 VDD.n5530 VSUBS 0.0867f
C12698 VDD.n5531 VSUBS 0.0867f
C12699 VDD.n5532 VSUBS 0.0867f
C12700 VDD.n5533 VSUBS 0.0867f
C12701 VDD.n5534 VSUBS 0.0867f
C12702 VDD.n5535 VSUBS 0.0867f
C12703 VDD.n5536 VSUBS 0.0867f
C12704 VDD.n5537 VSUBS 0.00723f
C12705 VDD.n5538 VSUBS 0.00354f
C12706 VDD.n5539 VSUBS 0.0145f
C12707 VDD.t128 VSUBS 0.0114f
C12708 VDD.t25 VSUBS 0.0114f
C12709 VDD.n5540 VSUBS 0.0268f
C12710 VDD.n5541 VSUBS 0.0126f
C12711 VDD.n5542 VSUBS 0.0264f
C12712 VDD.n5543 VSUBS 0.0142f
C12713 VDD.n5544 VSUBS 0.00723f
C12714 VDD.n5545 VSUBS 0.00354f
C12715 VDD.n5546 VSUBS 0.0145f
C12716 VDD.t77 VSUBS 0.0114f
C12717 VDD.t422 VSUBS 0.0114f
C12718 VDD.n5547 VSUBS 0.0268f
C12719 VDD.n5548 VSUBS 0.0126f
C12720 VDD.n5549 VSUBS 0.0264f
C12721 VDD.n5550 VSUBS 0.0142f
C12722 VDD.n5551 VSUBS 0.00723f
C12723 VDD.n5552 VSUBS 0.00354f
C12724 VDD.n5553 VSUBS 0.0145f
C12725 VDD.t84 VSUBS 0.0114f
C12726 VDD.t163 VSUBS 0.0114f
C12727 VDD.n5554 VSUBS 0.0268f
C12728 VDD.n5555 VSUBS 0.0126f
C12729 VDD.n5556 VSUBS 0.0264f
C12730 VDD.n5557 VSUBS 0.0142f
C12731 VDD.n5558 VSUBS 0.00723f
C12732 VDD.n5559 VSUBS 0.00354f
C12733 VDD.n5560 VSUBS 0.0145f
C12734 VDD.t74 VSUBS 0.0114f
C12735 VDD.t412 VSUBS 0.0114f
C12736 VDD.n5561 VSUBS 0.0268f
C12737 VDD.n5562 VSUBS 0.0126f
C12738 VDD.n5563 VSUBS 0.0264f
C12739 VDD.n5564 VSUBS 0.0142f
C12740 VDD.n5565 VSUBS 0.00723f
C12741 VDD.n5566 VSUBS 0.00354f
C12742 VDD.n5567 VSUBS 0.0145f
C12743 VDD.t109 VSUBS 0.0114f
C12744 VDD.t415 VSUBS 0.0114f
C12745 VDD.n5568 VSUBS 0.0268f
C12746 VDD.n5569 VSUBS 0.0126f
C12747 VDD.n5570 VSUBS 0.0264f
C12748 VDD.n5571 VSUBS 0.0142f
C12749 VDD.n5572 VSUBS 0.00723f
C12750 VDD.n5573 VSUBS 0.00354f
C12751 VDD.n5574 VSUBS 0.0145f
C12752 VDD.t399 VSUBS 0.0114f
C12753 VDD.t96 VSUBS 0.0114f
C12754 VDD.n5575 VSUBS 0.0268f
C12755 VDD.n5576 VSUBS 0.0126f
C12756 VDD.n5577 VSUBS 0.0264f
C12757 VDD.n5578 VSUBS 0.0142f
C12758 VDD.n5579 VSUBS 0.00723f
C12759 VDD.n5580 VSUBS 0.00354f
C12760 VDD.n5581 VSUBS 0.0145f
C12761 VDD.t395 VSUBS 0.0114f
C12762 VDD.t95 VSUBS 0.0114f
C12763 VDD.n5582 VSUBS 0.0268f
C12764 VDD.n5583 VSUBS 0.0126f
C12765 VDD.n5584 VSUBS 0.0264f
C12766 VDD.n5585 VSUBS 0.0142f
C12767 VDD.n5586 VSUBS 0.00723f
C12768 VDD.n5587 VSUBS 0.00354f
C12769 VDD.n5588 VSUBS 0.0145f
C12770 VDD.t75 VSUBS 0.0114f
C12771 VDD.t431 VSUBS 0.0114f
C12772 VDD.n5589 VSUBS 0.0268f
C12773 VDD.n5590 VSUBS 0.0126f
C12774 VDD.n5591 VSUBS 0.0264f
C12775 VDD.n5592 VSUBS 0.0142f
C12776 VDD.n5593 VSUBS 0.00723f
C12777 VDD.n5594 VSUBS 0.00354f
C12778 VDD.n5595 VSUBS 0.0145f
C12779 VDD.t455 VSUBS 0.0114f
C12780 VDD.t28 VSUBS 0.0114f
C12781 VDD.n5596 VSUBS 0.0268f
C12782 VDD.n5597 VSUBS 0.0126f
C12783 VDD.n5598 VSUBS 0.0264f
C12784 VDD.n5599 VSUBS 0.0142f
C12785 VDD.n5600 VSUBS 0.00723f
C12786 VDD.n5601 VSUBS 0.00354f
C12787 VDD.n5602 VSUBS 0.0145f
C12788 VDD.t26 VSUBS 0.0114f
C12789 VDD.t417 VSUBS 0.0114f
C12790 VDD.n5603 VSUBS 0.0268f
C12791 VDD.n5604 VSUBS 0.0126f
C12792 VDD.n5605 VSUBS 0.0264f
C12793 VDD.n5606 VSUBS 0.0142f
C12794 VDD.n5607 VSUBS 0.00723f
C12795 VDD.n5608 VSUBS 0.00354f
C12796 VDD.n5609 VSUBS 0.0145f
C12797 VDD.t34 VSUBS 0.0114f
C12798 VDD.t375 VSUBS 0.0114f
C12799 VDD.n5610 VSUBS 0.0268f
C12800 VDD.n5611 VSUBS 0.0126f
C12801 VDD.n5612 VSUBS 0.0264f
C12802 VDD.n5613 VSUBS 0.0142f
C12803 VDD.n5614 VSUBS 0.00723f
C12804 VDD.n5615 VSUBS 0.00354f
C12805 VDD.n5616 VSUBS 0.0145f
C12806 VDD.t451 VSUBS 0.0114f
C12807 VDD.t370 VSUBS 0.0114f
C12808 VDD.n5617 VSUBS 0.0268f
C12809 VDD.n5618 VSUBS 0.0126f
C12810 VDD.n5619 VSUBS 0.0264f
C12811 VDD.n5620 VSUBS 0.0142f
C12812 VDD.n5621 VSUBS 0.00723f
C12813 VDD.n5622 VSUBS 0.00354f
C12814 VDD.n5623 VSUBS 0.0145f
C12815 VDD.t404 VSUBS 0.0114f
C12816 VDD.t49 VSUBS 0.0114f
C12817 VDD.n5624 VSUBS 0.0268f
C12818 VDD.n5625 VSUBS 0.0126f
C12819 VDD.n5626 VSUBS 0.0264f
C12820 VDD.n5627 VSUBS 0.0142f
C12821 VDD.n5628 VSUBS 0.00723f
C12822 VDD.n5629 VSUBS 0.00354f
C12823 VDD.n5630 VSUBS 0.0145f
C12824 VDD.t92 VSUBS 0.0114f
C12825 VDD.t12 VSUBS 0.0114f
C12826 VDD.n5631 VSUBS 0.0268f
C12827 VDD.n5632 VSUBS 0.0126f
C12828 VDD.n5633 VSUBS 0.0264f
C12829 VDD.n5634 VSUBS 0.0142f
C12830 VDD.n5635 VSUBS 0.00723f
C12831 VDD.n5636 VSUBS 0.00354f
C12832 VDD.n5637 VSUBS 0.0145f
C12833 VDD.t41 VSUBS 0.0114f
C12834 VDD.t138 VSUBS 0.0114f
C12835 VDD.n5638 VSUBS 0.0268f
C12836 VDD.n5639 VSUBS 0.0126f
C12837 VDD.n5640 VSUBS 0.0264f
C12838 VDD.n5641 VSUBS 0.0142f
C12839 VDD.n5642 VSUBS 0.00723f
C12840 VDD.n5643 VSUBS 0.00354f
C12841 VDD.n5644 VSUBS 0.0145f
C12842 VDD.t86 VSUBS 0.0114f
C12843 VDD.t5 VSUBS 0.0114f
C12844 VDD.n5645 VSUBS 0.0268f
C12845 VDD.n5646 VSUBS 0.0126f
C12846 VDD.n5647 VSUBS 0.0264f
C12847 VDD.n5648 VSUBS 0.0142f
C12848 VDD.n5649 VSUBS 0.00723f
C12849 VDD.n5650 VSUBS 0.00354f
C12850 VDD.n5651 VSUBS 0.0145f
C12851 VDD.t425 VSUBS 0.0114f
C12852 VDD.t144 VSUBS 0.0114f
C12853 VDD.n5652 VSUBS 0.0268f
C12854 VDD.n5653 VSUBS 0.0126f
C12855 VDD.n5654 VSUBS 0.0264f
C12856 VDD.n5655 VSUBS 0.0142f
C12857 VDD.n5656 VSUBS 0.00723f
C12858 VDD.n5657 VSUBS 0.00354f
C12859 VDD.n5658 VSUBS 0.0145f
C12860 VDD.t386 VSUBS 0.0114f
C12861 VDD.t442 VSUBS 0.0114f
C12862 VDD.n5659 VSUBS 0.0268f
C12863 VDD.n5660 VSUBS 0.0126f
C12864 VDD.n5661 VSUBS 0.0264f
C12865 VDD.n5662 VSUBS 0.0142f
C12866 VDD.n5663 VSUBS 0.00723f
C12867 VDD.n5664 VSUBS 0.00354f
C12868 VDD.n5665 VSUBS 0.0145f
C12869 VDD.t44 VSUBS 0.0114f
C12870 VDD.t146 VSUBS 0.0114f
C12871 VDD.n5666 VSUBS 0.0268f
C12872 VDD.n5667 VSUBS 0.0126f
C12873 VDD.n5668 VSUBS 0.0264f
C12874 VDD.n5669 VSUBS 0.0142f
C12875 VDD.n5670 VSUBS 0.00723f
C12876 VDD.n5671 VSUBS 0.00354f
C12877 VDD.n5672 VSUBS 0.0202f
C12878 VDD.t430 VSUBS 0.0114f
C12879 VDD.t440 VSUBS 0.0114f
C12880 VDD.n5673 VSUBS 0.0268f
C12881 VDD.n5674 VSUBS 0.0126f
C12882 VDD.n5675 VSUBS 0.0264f
C12883 VDD.n5676 VSUBS 0.0142f
C12884 VDD.n5677 VSUBS 0.215f
C12885 VDD.n5678 VSUBS 0.0867f
C12886 VDD.n5679 VSUBS 0.0867f
C12887 VDD.n5680 VSUBS 0.0867f
C12888 VDD.n5681 VSUBS 0.0867f
C12889 VDD.n5682 VSUBS 0.0867f
C12890 VDD.n5683 VSUBS 0.0867f
C12891 VDD.n5684 VSUBS 0.0867f
C12892 VDD.n5685 VSUBS 0.0867f
C12893 VDD.n5686 VSUBS 0.0867f
C12894 VDD.n5687 VSUBS 0.0867f
C12895 VDD.n5688 VSUBS 0.0867f
C12896 VDD.n5689 VSUBS 0.0867f
C12897 VDD.n5690 VSUBS 0.0867f
C12898 VDD.n5691 VSUBS 0.0867f
C12899 VDD.n5692 VSUBS 0.0867f
C12900 VDD.n5693 VSUBS 0.0867f
C12901 VDD.n5694 VSUBS 0.0867f
C12902 VDD.n5695 VSUBS 0.0867f
C12903 VDD.n5696 VSUBS 0.0867f
C12904 VDD.n5697 VSUBS 0.0867f
C12905 VDD.n5698 VSUBS 0.0867f
C12906 VDD.n5699 VSUBS 0.0867f
C12907 VDD.n5700 VSUBS 0.0867f
C12908 VDD.n5701 VSUBS 0.0867f
C12909 VDD.n5702 VSUBS 0.0867f
C12910 VDD.n5703 VSUBS 0.0867f
C12911 VDD.n5704 VSUBS 0.0867f
C12912 VDD.n5705 VSUBS 0.0867f
C12913 VDD.n5706 VSUBS 0.0867f
C12914 VDD.n5707 VSUBS 0.0867f
C12915 VDD.n5708 VSUBS 0.0867f
C12916 VDD.n5709 VSUBS 0.0867f
C12917 VDD.n5710 VSUBS 0.0867f
C12918 VDD.n5711 VSUBS 0.0867f
C12919 VDD.n5712 VSUBS 0.0867f
C12920 VDD.n5713 VSUBS 0.0867f
C12921 VDD.n5714 VSUBS 0.0867f
C12922 VDD.n5715 VSUBS 0.0867f
C12923 VDD.n5716 VSUBS 0.00723f
C12924 VDD.n5717 VSUBS 0.00354f
C12925 VDD.n5718 VSUBS 0.0145f
C12926 VDD.t441 VSUBS 0.0114f
C12927 VDD.t108 VSUBS 0.0114f
C12928 VDD.n5719 VSUBS 0.0268f
C12929 VDD.n5720 VSUBS 0.0127f
C12930 VDD.n5721 VSUBS 0.0267f
C12931 VDD.n5722 VSUBS 0.0142f
C12932 VDD.n5723 VSUBS 0.00723f
C12933 VDD.n5724 VSUBS 0.00354f
C12934 VDD.n5725 VSUBS 0.0145f
C12935 VDD.t418 VSUBS 0.0114f
C12936 VDD.t118 VSUBS 0.0114f
C12937 VDD.n5726 VSUBS 0.0268f
C12938 VDD.n5727 VSUBS 0.0127f
C12939 VDD.n5728 VSUBS 0.0267f
C12940 VDD.n5729 VSUBS 0.0142f
C12941 VDD.n5730 VSUBS 0.00723f
C12942 VDD.n5731 VSUBS 0.00354f
C12943 VDD.n5732 VSUBS 0.0145f
C12944 VDD.t164 VSUBS 0.0114f
C12945 VDD.t382 VSUBS 0.0114f
C12946 VDD.n5733 VSUBS 0.0268f
C12947 VDD.n5734 VSUBS 0.0127f
C12948 VDD.n5735 VSUBS 0.0267f
C12949 VDD.n5736 VSUBS 0.0142f
C12950 VDD.n5737 VSUBS 0.00723f
C12951 VDD.n5738 VSUBS 0.00354f
C12952 VDD.n5739 VSUBS 0.0145f
C12953 VDD.t406 VSUBS 0.0114f
C12954 VDD.t388 VSUBS 0.0114f
C12955 VDD.n5740 VSUBS 0.0268f
C12956 VDD.n5741 VSUBS 0.0127f
C12957 VDD.n5742 VSUBS 0.0267f
C12958 VDD.n5743 VSUBS 0.0142f
C12959 VDD.n5744 VSUBS 0.00723f
C12960 VDD.n5745 VSUBS 0.00354f
C12961 VDD.n5746 VSUBS 0.0145f
C12962 VDD.t437 VSUBS 0.0114f
C12963 VDD.t112 VSUBS 0.0114f
C12964 VDD.n5747 VSUBS 0.0268f
C12965 VDD.n5748 VSUBS 0.0127f
C12966 VDD.n5749 VSUBS 0.0267f
C12967 VDD.n5750 VSUBS 0.0142f
C12968 VDD.n5751 VSUBS 0.00723f
C12969 VDD.n5752 VSUBS 0.00354f
C12970 VDD.n5753 VSUBS 0.0145f
C12971 VDD.t116 VSUBS 0.0114f
C12972 VDD.t114 VSUBS 0.0114f
C12973 VDD.n5754 VSUBS 0.0268f
C12974 VDD.n5755 VSUBS 0.0127f
C12975 VDD.n5756 VSUBS 0.0267f
C12976 VDD.n5757 VSUBS 0.0142f
C12977 VDD.n5758 VSUBS 0.00723f
C12978 VDD.n5759 VSUBS 0.00354f
C12979 VDD.n5760 VSUBS 0.0145f
C12980 VDD.t66 VSUBS 0.0114f
C12981 VDD.t148 VSUBS 0.0114f
C12982 VDD.n5761 VSUBS 0.0268f
C12983 VDD.n5762 VSUBS 0.0127f
C12984 VDD.n5763 VSUBS 0.0267f
C12985 VDD.n5764 VSUBS 0.0142f
C12986 VDD.n5765 VSUBS 0.00723f
C12987 VDD.n5766 VSUBS 0.00354f
C12988 VDD.n5767 VSUBS 0.0145f
C12989 VDD.t434 VSUBS 0.0114f
C12990 VDD.t123 VSUBS 0.0114f
C12991 VDD.n5768 VSUBS 0.0268f
C12992 VDD.n5769 VSUBS 0.0127f
C12993 VDD.n5770 VSUBS 0.0267f
C12994 VDD.n5771 VSUBS 0.0142f
C12995 VDD.n5772 VSUBS 0.00723f
C12996 VDD.n5773 VSUBS 0.00354f
C12997 VDD.n5774 VSUBS 0.0145f
C12998 VDD.t102 VSUBS 0.0114f
C12999 VDD.t409 VSUBS 0.0114f
C13000 VDD.n5775 VSUBS 0.0268f
C13001 VDD.n5776 VSUBS 0.0127f
C13002 VDD.n5777 VSUBS 0.0267f
C13003 VDD.n5778 VSUBS 0.0142f
C13004 VDD.n5779 VSUBS 0.00723f
C13005 VDD.n5780 VSUBS 0.00354f
C13006 VDD.n5781 VSUBS 0.0145f
C13007 VDD.t416 VSUBS 0.0114f
C13008 VDD.t130 VSUBS 0.0114f
C13009 VDD.n5782 VSUBS 0.0268f
C13010 VDD.n5783 VSUBS 0.0127f
C13011 VDD.n5784 VSUBS 0.0267f
C13012 VDD.n5785 VSUBS 0.0142f
C13013 VDD.n5786 VSUBS 0.00723f
C13014 VDD.n5787 VSUBS 0.00354f
C13015 VDD.n5788 VSUBS 0.0145f
C13016 VDD.t119 VSUBS 0.0114f
C13017 VDD.t147 VSUBS 0.0114f
C13018 VDD.n5789 VSUBS 0.0268f
C13019 VDD.n5790 VSUBS 0.0127f
C13020 VDD.n5791 VSUBS 0.0267f
C13021 VDD.n5792 VSUBS 0.0142f
C13022 VDD.n5793 VSUBS 0.00723f
C13023 VDD.n5794 VSUBS 0.00354f
C13024 VDD.n5795 VSUBS 0.0145f
C13025 VDD.t445 VSUBS 0.0114f
C13026 VDD.t421 VSUBS 0.0114f
C13027 VDD.n5796 VSUBS 0.0268f
C13028 VDD.n5797 VSUBS 0.0127f
C13029 VDD.n5798 VSUBS 0.0267f
C13030 VDD.n5799 VSUBS 0.0142f
C13031 VDD.n5800 VSUBS 0.00723f
C13032 VDD.n5801 VSUBS 0.00354f
C13033 VDD.n5802 VSUBS 0.0145f
C13034 VDD.t374 VSUBS 0.0114f
C13035 VDD.t65 VSUBS 0.0114f
C13036 VDD.n5803 VSUBS 0.0268f
C13037 VDD.n5804 VSUBS 0.0127f
C13038 VDD.n5805 VSUBS 0.0267f
C13039 VDD.n5806 VSUBS 0.0142f
C13040 VDD.n5807 VSUBS 0.00723f
C13041 VDD.n5808 VSUBS 0.00354f
C13042 VDD.n5809 VSUBS 0.0145f
C13043 VDD.t113 VSUBS 0.0114f
C13044 VDD.t126 VSUBS 0.0114f
C13045 VDD.n5810 VSUBS 0.0268f
C13046 VDD.n5811 VSUBS 0.0127f
C13047 VDD.n5812 VSUBS 0.0267f
C13048 VDD.n5813 VSUBS 0.0142f
C13049 VDD.n5814 VSUBS 0.00723f
C13050 VDD.n5815 VSUBS 0.00354f
C13051 VDD.n5816 VSUBS 0.0145f
C13052 VDD.t67 VSUBS 0.0114f
C13053 VDD.t429 VSUBS 0.0114f
C13054 VDD.n5817 VSUBS 0.0268f
C13055 VDD.n5818 VSUBS 0.0127f
C13056 VDD.n5819 VSUBS 0.0267f
C13057 VDD.n5820 VSUBS 0.0142f
C13058 VDD.n5821 VSUBS 0.00723f
C13059 VDD.n5822 VSUBS 0.00354f
C13060 VDD.n5823 VSUBS 0.0145f
C13061 VDD.t401 VSUBS 0.0114f
C13062 VDD.t64 VSUBS 0.0114f
C13063 VDD.n5824 VSUBS 0.0268f
C13064 VDD.n5825 VSUBS 0.0127f
C13065 VDD.n5826 VSUBS 0.0267f
C13066 VDD.n5827 VSUBS 0.0142f
C13067 VDD.n5828 VSUBS 0.00723f
C13068 VDD.n5829 VSUBS 0.00354f
C13069 VDD.n5830 VSUBS 0.0145f
C13070 VDD.t373 VSUBS 0.0114f
C13071 VDD.t407 VSUBS 0.0114f
C13072 VDD.n5831 VSUBS 0.0268f
C13073 VDD.n5832 VSUBS 0.0127f
C13074 VDD.n5833 VSUBS 0.0267f
C13075 VDD.n5834 VSUBS 0.0142f
C13076 VDD.n5835 VSUBS 0.00723f
C13077 VDD.n5836 VSUBS 0.00354f
C13078 VDD.n5837 VSUBS 0.0145f
C13079 VDD.t132 VSUBS 0.0114f
C13080 VDD.t30 VSUBS 0.0114f
C13081 VDD.n5838 VSUBS 0.0268f
C13082 VDD.n5839 VSUBS 0.0127f
C13083 VDD.n5840 VSUBS 0.0267f
C13084 VDD.n5841 VSUBS 0.0142f
C13085 VDD.n5842 VSUBS 0.00723f
C13086 VDD.n5843 VSUBS 0.00354f
C13087 VDD.n5844 VSUBS 0.0145f
C13088 VDD.t403 VSUBS 0.0114f
C13089 VDD.t46 VSUBS 0.0114f
C13090 VDD.n5845 VSUBS 0.0268f
C13091 VDD.n5846 VSUBS 0.0127f
C13092 VDD.n5847 VSUBS 0.0267f
C13093 VDD.n5848 VSUBS 0.0142f
C13094 VDD.n5849 VSUBS 0.00723f
C13095 VDD.n5850 VSUBS 0.00354f
C13096 VDD.n5851 VSUBS 0.0202f
C13097 VDD.t402 VSUBS 0.0114f
C13098 VDD.t448 VSUBS 0.0114f
C13099 VDD.n5852 VSUBS 0.0268f
C13100 VDD.n5853 VSUBS 0.0127f
C13101 VDD.n5854 VSUBS 0.0267f
C13102 VDD.n5855 VSUBS 0.0142f
C13103 VDD.n5856 VSUBS 0.215f
C13104 VDD.n5857 VSUBS 0.0867f
C13105 VDD.n5858 VSUBS 0.0867f
C13106 VDD.n5859 VSUBS 0.0867f
C13107 VDD.n5860 VSUBS 0.0867f
C13108 VDD.n5861 VSUBS 0.0867f
C13109 VDD.n5862 VSUBS 0.0867f
C13110 VDD.n5863 VSUBS 0.0867f
C13111 VDD.n5864 VSUBS 0.0867f
C13112 VDD.n5865 VSUBS 0.0867f
C13113 VDD.n5866 VSUBS 0.0867f
C13114 VDD.n5867 VSUBS 0.0867f
C13115 VDD.n5868 VSUBS 0.0867f
C13116 VDD.n5869 VSUBS 0.0867f
C13117 VDD.n5870 VSUBS 0.0867f
C13118 VDD.n5871 VSUBS 0.0867f
C13119 VDD.n5872 VSUBS 0.0867f
C13120 VDD.n5873 VSUBS 0.0867f
C13121 VDD.n5874 VSUBS 0.0867f
C13122 VDD.n5875 VSUBS 0.0867f
C13123 VDD.n5876 VSUBS 0.0867f
C13124 VDD.n5877 VSUBS 0.0867f
C13125 VDD.n5878 VSUBS 0.0867f
C13126 VDD.n5879 VSUBS 0.0867f
C13127 VDD.n5880 VSUBS 0.0867f
C13128 VDD.n5881 VSUBS 0.0867f
C13129 VDD.n5882 VSUBS 0.0867f
C13130 VDD.n5883 VSUBS 0.0867f
C13131 VDD.n5884 VSUBS 0.0867f
C13132 VDD.n5885 VSUBS 0.0867f
C13133 VDD.n5886 VSUBS 0.0867f
C13134 VDD.n5887 VSUBS 0.0867f
C13135 VDD.n5888 VSUBS 0.0867f
C13136 VDD.n5889 VSUBS 0.0867f
C13137 VDD.n5890 VSUBS 0.0867f
C13138 VDD.n5891 VSUBS 0.0867f
C13139 VDD.n5892 VSUBS 0.0867f
C13140 VDD.n5893 VSUBS 0.0867f
C13141 VDD.n5894 VSUBS 0.0867f
C13142 VDD.n5895 VSUBS 0.00737f
C13143 VDD.n5896 VSUBS 0.00365f
C13144 VDD.n5897 VSUBS 0.0145f
C13145 VDD.t447 VSUBS 0.0114f
C13146 VDD.t32 VSUBS 0.0114f
C13147 VDD.n5898 VSUBS 0.0268f
C13148 VDD.n5899 VSUBS 0.0123f
C13149 VDD.n5900 VSUBS 0.0254f
C13150 VDD.n5901 VSUBS 0.0142f
C13151 VDD.n5902 VSUBS 0.00737f
C13152 VDD.n5903 VSUBS 0.00365f
C13153 VDD.n5904 VSUBS 0.0145f
C13154 VDD.t392 VSUBS 0.0114f
C13155 VDD.t125 VSUBS 0.0114f
C13156 VDD.n5905 VSUBS 0.0268f
C13157 VDD.n5906 VSUBS 0.0123f
C13158 VDD.n5907 VSUBS 0.0254f
C13159 VDD.n5908 VSUBS 0.0142f
C13160 VDD.n5909 VSUBS 0.00737f
C13161 VDD.n5910 VSUBS 0.00365f
C13162 VDD.n5911 VSUBS 0.0145f
C13163 VDD.t438 VSUBS 0.0114f
C13164 VDD.t457 VSUBS 0.0114f
C13165 VDD.n5912 VSUBS 0.0268f
C13166 VDD.n5913 VSUBS 0.0123f
C13167 VDD.n5914 VSUBS 0.0254f
C13168 VDD.n5915 VSUBS 0.0142f
C13169 VDD.n5916 VSUBS 0.00737f
C13170 VDD.n5917 VSUBS 0.00365f
C13171 VDD.n5918 VSUBS 0.0145f
C13172 VDD.t454 VSUBS 0.0114f
C13173 VDD.t420 VSUBS 0.0114f
C13174 VDD.n5919 VSUBS 0.0268f
C13175 VDD.n5920 VSUBS 0.0123f
C13176 VDD.n5921 VSUBS 0.0254f
C13177 VDD.n5922 VSUBS 0.0142f
C13178 VDD.n5923 VSUBS 0.00737f
C13179 VDD.n5924 VSUBS 0.00365f
C13180 VDD.n5925 VSUBS 0.0145f
C13181 VDD.t379 VSUBS 0.0114f
C13182 VDD.t426 VSUBS 0.0114f
C13183 VDD.n5926 VSUBS 0.0268f
C13184 VDD.n5927 VSUBS 0.0123f
C13185 VDD.n5928 VSUBS 0.0254f
C13186 VDD.n5929 VSUBS 0.0142f
C13187 VDD.n5930 VSUBS 0.00737f
C13188 VDD.n5931 VSUBS 0.00365f
C13189 VDD.n5932 VSUBS 0.0145f
C13190 VDD.t377 VSUBS 0.0114f
C13191 VDD.t94 VSUBS 0.0114f
C13192 VDD.n5933 VSUBS 0.0268f
C13193 VDD.n5934 VSUBS 0.0123f
C13194 VDD.n5935 VSUBS 0.0254f
C13195 VDD.n5936 VSUBS 0.0142f
C13196 VDD.n5937 VSUBS 0.00737f
C13197 VDD.n5938 VSUBS 0.00365f
C13198 VDD.n5939 VSUBS 0.0145f
C13199 VDD.t51 VSUBS 0.0114f
C13200 VDD.t427 VSUBS 0.0114f
C13201 VDD.n5940 VSUBS 0.0268f
C13202 VDD.n5941 VSUBS 0.0123f
C13203 VDD.n5942 VSUBS 0.0254f
C13204 VDD.n5943 VSUBS 0.0142f
C13205 VDD.n5944 VSUBS 0.00737f
C13206 VDD.n5945 VSUBS 0.00365f
C13207 VDD.n5946 VSUBS 0.0145f
C13208 VDD.t390 VSUBS 0.0114f
C13209 VDD.t111 VSUBS 0.0114f
C13210 VDD.n5947 VSUBS 0.0268f
C13211 VDD.n5948 VSUBS 0.0123f
C13212 VDD.n5949 VSUBS 0.0254f
C13213 VDD.n5950 VSUBS 0.0142f
C13214 VDD.n5951 VSUBS 0.00737f
C13215 VDD.n5952 VSUBS 0.00365f
C13216 VDD.n5953 VSUBS 0.0145f
C13217 VDD.t85 VSUBS 0.0114f
C13218 VDD.t90 VSUBS 0.0114f
C13219 VDD.n5954 VSUBS 0.0268f
C13220 VDD.n5955 VSUBS 0.0123f
C13221 VDD.n5956 VSUBS 0.0254f
C13222 VDD.n5957 VSUBS 0.0142f
C13223 VDD.n5958 VSUBS 0.00737f
C13224 VDD.n5959 VSUBS 0.00365f
C13225 VDD.n5960 VSUBS 0.0145f
C13226 VDD.t145 VSUBS 0.0114f
C13227 VDD.t154 VSUBS 0.0114f
C13228 VDD.n5961 VSUBS 0.0268f
C13229 VDD.n5962 VSUBS 0.0123f
C13230 VDD.n5963 VSUBS 0.0254f
C13231 VDD.n5964 VSUBS 0.0142f
C13232 VDD.n5965 VSUBS 0.00737f
C13233 VDD.n5966 VSUBS 0.00365f
C13234 VDD.n5967 VSUBS 0.0145f
C13235 VDD.t69 VSUBS 0.0114f
C13236 VDD.t106 VSUBS 0.0114f
C13237 VDD.n5968 VSUBS 0.0268f
C13238 VDD.n5969 VSUBS 0.0123f
C13239 VDD.n5970 VSUBS 0.0254f
C13240 VDD.n5971 VSUBS 0.0142f
C13241 VDD.n5972 VSUBS 0.00737f
C13242 VDD.n5973 VSUBS 0.00365f
C13243 VDD.n5974 VSUBS 0.0145f
C13244 VDD.t150 VSUBS 0.0114f
C13245 VDD.t134 VSUBS 0.0114f
C13246 VDD.n5975 VSUBS 0.0268f
C13247 VDD.n5976 VSUBS 0.0123f
C13248 VDD.n5977 VSUBS 0.0254f
C13249 VDD.n5978 VSUBS 0.0142f
C13250 VDD.n5979 VSUBS 0.00737f
C13251 VDD.n5980 VSUBS 0.00365f
C13252 VDD.n5981 VSUBS 0.0145f
C13253 VDD.t439 VSUBS 0.0114f
C13254 VDD.t433 VSUBS 0.0114f
C13255 VDD.n5982 VSUBS 0.0268f
C13256 VDD.n5983 VSUBS 0.0123f
C13257 VDD.n5984 VSUBS 0.0254f
C13258 VDD.n5985 VSUBS 0.0142f
C13259 VDD.n5986 VSUBS 0.00737f
C13260 VDD.n5987 VSUBS 0.00365f
C13261 VDD.n5988 VSUBS 0.0145f
C13262 VDD.t166 VSUBS 0.0114f
C13263 VDD.t410 VSUBS 0.0114f
C13264 VDD.n5989 VSUBS 0.0268f
C13265 VDD.n5990 VSUBS 0.0123f
C13266 VDD.n5991 VSUBS 0.0254f
C13267 VDD.n5992 VSUBS 0.0142f
C13268 VDD.n5993 VSUBS 0.00737f
C13269 VDD.n5994 VSUBS 0.00365f
C13270 VDD.n5995 VSUBS 0.0145f
C13271 VDD.t1 VSUBS 0.0114f
C13272 VDD.t453 VSUBS 0.0114f
C13273 VDD.n5996 VSUBS 0.0268f
C13274 VDD.n5997 VSUBS 0.0123f
C13275 VDD.n5998 VSUBS 0.0254f
C13276 VDD.n5999 VSUBS 0.0142f
C13277 VDD.n6000 VSUBS 0.00737f
C13278 VDD.n6001 VSUBS 0.00365f
C13279 VDD.n6002 VSUBS 0.0145f
C13280 VDD.t124 VSUBS 0.0114f
C13281 VDD.t432 VSUBS 0.0114f
C13282 VDD.n6003 VSUBS 0.0268f
C13283 VDD.n6004 VSUBS 0.0123f
C13284 VDD.n6005 VSUBS 0.0254f
C13285 VDD.n6006 VSUBS 0.0142f
C13286 VDD.n6007 VSUBS 0.00737f
C13287 VDD.n6008 VSUBS 0.00365f
C13288 VDD.n6009 VSUBS 0.0145f
C13289 VDD.t369 VSUBS 0.0114f
C13290 VDD.t149 VSUBS 0.0114f
C13291 VDD.n6010 VSUBS 0.0268f
C13292 VDD.n6011 VSUBS 0.0123f
C13293 VDD.n6012 VSUBS 0.0254f
C13294 VDD.n6013 VSUBS 0.0142f
C13295 VDD.n6014 VSUBS 0.00737f
C13296 VDD.n6015 VSUBS 0.00365f
C13297 VDD.n6016 VSUBS 0.0145f
C13298 VDD.t89 VSUBS 0.0114f
C13299 VDD.t396 VSUBS 0.0114f
C13300 VDD.n6017 VSUBS 0.0268f
C13301 VDD.n6018 VSUBS 0.0123f
C13302 VDD.n6019 VSUBS 0.0254f
C13303 VDD.n6020 VSUBS 0.0142f
C13304 VDD.n6021 VSUBS 0.00737f
C13305 VDD.n6022 VSUBS 0.00365f
C13306 VDD.n6023 VSUBS 0.0145f
C13307 VDD.t400 VSUBS 0.0114f
C13308 VDD.t103 VSUBS 0.0114f
C13309 VDD.n6024 VSUBS 0.0268f
C13310 VDD.n6025 VSUBS 0.0123f
C13311 VDD.n6026 VSUBS 0.0254f
C13312 VDD.n6027 VSUBS 0.0142f
C13313 VDD.n6028 VSUBS 0.00737f
C13314 VDD.n6029 VSUBS 0.00365f
C13315 VDD.n6030 VSUBS 0.0202f
C13316 VDD.t424 VSUBS 0.0114f
C13317 VDD.t62 VSUBS 0.0114f
C13318 VDD.n6031 VSUBS 0.0268f
C13319 VDD.n6032 VSUBS 0.0123f
C13320 VDD.n6033 VSUBS 0.0254f
C13321 VDD.n6034 VSUBS 0.0142f
C13322 VDD.n6035 VSUBS 0.215f
C13323 VDD.n6036 VSUBS 0.0867f
C13324 VDD.n6037 VSUBS 0.0867f
C13325 VDD.n6038 VSUBS 0.0867f
C13326 VDD.n6039 VSUBS 0.0867f
C13327 VDD.n6040 VSUBS 0.0867f
C13328 VDD.n6041 VSUBS 0.0867f
C13329 VDD.n6042 VSUBS 0.0867f
C13330 VDD.n6043 VSUBS 0.0867f
C13331 VDD.n6044 VSUBS 0.0867f
C13332 VDD.n6045 VSUBS 0.0867f
C13333 VDD.n6046 VSUBS 0.0867f
C13334 VDD.n6047 VSUBS 0.0867f
C13335 VDD.n6048 VSUBS 0.0867f
C13336 VDD.n6049 VSUBS 0.0867f
C13337 VDD.n6050 VSUBS 0.0867f
C13338 VDD.n6051 VSUBS 0.0867f
C13339 VDD.n6052 VSUBS 0.0867f
C13340 VDD.n6053 VSUBS 0.0867f
C13341 VDD.n6054 VSUBS 0.0867f
C13342 VDD.n6055 VSUBS 0.0867f
C13343 VDD.n6056 VSUBS 0.0867f
C13344 VDD.n6057 VSUBS 0.0867f
C13345 VDD.n6058 VSUBS 0.0867f
C13346 VDD.n6059 VSUBS 0.0867f
C13347 VDD.n6060 VSUBS 0.0867f
C13348 VDD.n6061 VSUBS 0.0867f
C13349 VDD.n6062 VSUBS 0.0867f
C13350 VDD.n6063 VSUBS 0.0867f
C13351 VDD.n6064 VSUBS 0.0867f
C13352 VDD.n6065 VSUBS 0.0867f
C13353 VDD.n6066 VSUBS 0.0867f
C13354 VDD.n6067 VSUBS 0.0867f
C13355 VDD.n6068 VSUBS 0.0867f
C13356 VDD.n6069 VSUBS 0.0867f
C13357 VDD.n6070 VSUBS 0.0867f
C13358 VDD.n6071 VSUBS 0.0867f
C13359 VDD.n6072 VSUBS 0.0867f
C13360 VDD.n6073 VSUBS 0.0867f
C13361 VDD.n6074 VSUBS 0.0075f
C13362 VDD.n6075 VSUBS 0.00379f
C13363 VDD.n6076 VSUBS 0.0145f
C13364 VDD.t121 VSUBS 0.0114f
C13365 VDD.t385 VSUBS 0.0114f
C13366 VDD.n6077 VSUBS 0.0268f
C13367 VDD.n6078 VSUBS 0.0118f
C13368 VDD.n6079 VSUBS 0.0242f
C13369 VDD.n6080 VSUBS 0.0142f
C13370 VDD.n6081 VSUBS 0.0075f
C13371 VDD.n6082 VSUBS 0.00379f
C13372 VDD.n6083 VSUBS 0.0145f
C13373 VDD.t459 VSUBS 0.0114f
C13374 VDD.t381 VSUBS 0.0114f
C13375 VDD.n6084 VSUBS 0.0268f
C13376 VDD.n6085 VSUBS 0.0118f
C13377 VDD.n6086 VSUBS 0.0242f
C13378 VDD.n6087 VSUBS 0.0142f
C13379 VDD.n6088 VSUBS 0.0075f
C13380 VDD.n6089 VSUBS 0.00379f
C13381 VDD.n6090 VSUBS 0.0145f
C13382 VDD.t104 VSUBS 0.0114f
C13383 VDD.t139 VSUBS 0.0114f
C13384 VDD.n6091 VSUBS 0.0268f
C13385 VDD.n6092 VSUBS 0.0118f
C13386 VDD.n6093 VSUBS 0.0242f
C13387 VDD.n6094 VSUBS 0.0142f
C13388 VDD.n6095 VSUBS 0.0075f
C13389 VDD.n6096 VSUBS 0.00379f
C13390 VDD.n6097 VSUBS 0.0145f
C13391 VDD.t3 VSUBS 0.0114f
C13392 VDD.t413 VSUBS 0.0114f
C13393 VDD.n6098 VSUBS 0.0268f
C13394 VDD.n6099 VSUBS 0.0118f
C13395 VDD.n6100 VSUBS 0.0242f
C13396 VDD.n6101 VSUBS 0.0142f
C13397 VDD.n6102 VSUBS 0.0075f
C13398 VDD.n6103 VSUBS 0.00379f
C13399 VDD.n6104 VSUBS 0.0145f
C13400 VDD.t16 VSUBS 0.0114f
C13401 VDD.t9 VSUBS 0.0114f
C13402 VDD.n6105 VSUBS 0.0268f
C13403 VDD.n6106 VSUBS 0.0118f
C13404 VDD.n6107 VSUBS 0.0242f
C13405 VDD.n6108 VSUBS 0.0142f
C13406 VDD.n6109 VSUBS 0.0075f
C13407 VDD.n6110 VSUBS 0.00379f
C13408 VDD.n6111 VSUBS 0.0145f
C13409 VDD.t387 VSUBS 0.0114f
C13410 VDD.t449 VSUBS 0.0114f
C13411 VDD.n6112 VSUBS 0.0268f
C13412 VDD.n6113 VSUBS 0.0118f
C13413 VDD.n6114 VSUBS 0.0242f
C13414 VDD.n6115 VSUBS 0.0142f
C13415 VDD.n6116 VSUBS 0.0075f
C13416 VDD.n6117 VSUBS 0.00379f
C13417 VDD.n6118 VSUBS 0.0145f
C13418 VDD.t372 VSUBS 0.0114f
C13419 VDD.t107 VSUBS 0.0114f
C13420 VDD.n6119 VSUBS 0.0268f
C13421 VDD.n6120 VSUBS 0.0118f
C13422 VDD.n6121 VSUBS 0.0242f
C13423 VDD.n6122 VSUBS 0.0142f
C13424 VDD.n6123 VSUBS 0.0075f
C13425 VDD.n6124 VSUBS 0.00379f
C13426 VDD.n6125 VSUBS 0.0145f
C13427 VDD.t97 VSUBS 0.0114f
C13428 VDD.t371 VSUBS 0.0114f
C13429 VDD.n6126 VSUBS 0.0268f
C13430 VDD.n6127 VSUBS 0.0118f
C13431 VDD.n6128 VSUBS 0.0242f
C13432 VDD.n6129 VSUBS 0.0142f
C13433 VDD.n6130 VSUBS 0.0075f
C13434 VDD.n6131 VSUBS 0.00379f
C13435 VDD.n6132 VSUBS 0.0145f
C13436 VDD.t122 VSUBS 0.0114f
C13437 VDD.t384 VSUBS 0.0114f
C13438 VDD.n6133 VSUBS 0.0268f
C13439 VDD.n6134 VSUBS 0.0118f
C13440 VDD.n6135 VSUBS 0.0242f
C13441 VDD.n6136 VSUBS 0.0142f
C13442 VDD.n6137 VSUBS 0.0075f
C13443 VDD.n6138 VSUBS 0.00379f
C13444 VDD.n6139 VSUBS 0.0145f
C13445 VDD.t393 VSUBS 0.0114f
C13446 VDD.t131 VSUBS 0.0114f
C13447 VDD.n6140 VSUBS 0.0268f
C13448 VDD.n6141 VSUBS 0.0118f
C13449 VDD.n6142 VSUBS 0.0242f
C13450 VDD.n6143 VSUBS 0.0142f
C13451 VDD.n6144 VSUBS 0.0075f
C13452 VDD.n6145 VSUBS 0.00379f
C13453 VDD.n6146 VSUBS 0.0145f
C13454 VDD.t464 VSUBS 0.0114f
C13455 VDD.t463 VSUBS 0.0114f
C13456 VDD.n6147 VSUBS 0.0268f
C13457 VDD.n6148 VSUBS 0.0118f
C13458 VDD.n6149 VSUBS 0.0242f
C13459 VDD.n6150 VSUBS 0.0142f
C13460 VDD.n6151 VSUBS 0.0075f
C13461 VDD.n6152 VSUBS 0.00379f
C13462 VDD.n6153 VSUBS 0.0145f
C13463 VDD.t136 VSUBS 0.0114f
C13464 VDD.t376 VSUBS 0.0114f
C13465 VDD.n6154 VSUBS 0.0268f
C13466 VDD.n6155 VSUBS 0.0118f
C13467 VDD.n6156 VSUBS 0.0242f
C13468 VDD.n6157 VSUBS 0.0142f
C13469 VDD.n6158 VSUBS 0.0075f
C13470 VDD.n6159 VSUBS 0.00379f
C13471 VDD.n6160 VSUBS 0.0145f
C13472 VDD.t73 VSUBS 0.0114f
C13473 VDD.t48 VSUBS 0.0114f
C13474 VDD.n6161 VSUBS 0.0268f
C13475 VDD.n6162 VSUBS 0.0118f
C13476 VDD.n6163 VSUBS 0.0242f
C13477 VDD.n6164 VSUBS 0.0142f
C13478 VDD.n6165 VSUBS 0.0075f
C13479 VDD.n6166 VSUBS 0.00379f
C13480 VDD.n6167 VSUBS 0.0145f
C13481 VDD.t137 VSUBS 0.0114f
C13482 VDD.t87 VSUBS 0.0114f
C13483 VDD.n6168 VSUBS 0.0268f
C13484 VDD.n6169 VSUBS 0.0118f
C13485 VDD.n6170 VSUBS 0.0242f
C13486 VDD.n6171 VSUBS 0.0142f
C13487 VDD.n6172 VSUBS 0.0075f
C13488 VDD.n6173 VSUBS 0.00379f
C13489 VDD.n6174 VSUBS 0.0145f
C13490 VDD.t10 VSUBS 0.0114f
C13491 VDD.t20 VSUBS 0.0114f
C13492 VDD.n6175 VSUBS 0.0268f
C13493 VDD.n6176 VSUBS 0.0118f
C13494 VDD.n6177 VSUBS 0.0242f
C13495 VDD.n6178 VSUBS 0.0142f
C13496 VDD.n6179 VSUBS 0.0075f
C13497 VDD.n6180 VSUBS 0.00379f
C13498 VDD.n6181 VSUBS 0.0145f
C13499 VDD.t398 VSUBS 0.0114f
C13500 VDD.t82 VSUBS 0.0114f
C13501 VDD.n6182 VSUBS 0.0268f
C13502 VDD.n6183 VSUBS 0.0118f
C13503 VDD.n6184 VSUBS 0.0242f
C13504 VDD.n6185 VSUBS 0.0142f
C13505 VDD.n6186 VSUBS 0.0075f
C13506 VDD.n6187 VSUBS 0.00379f
C13507 VDD.n6188 VSUBS 0.0145f
C13508 VDD.t383 VSUBS 0.0114f
C13509 VDD.t151 VSUBS 0.0114f
C13510 VDD.n6189 VSUBS 0.0268f
C13511 VDD.n6190 VSUBS 0.0118f
C13512 VDD.n6191 VSUBS 0.0242f
C13513 VDD.n6192 VSUBS 0.0142f
C13514 VDD.n6193 VSUBS 0.0075f
C13515 VDD.n6194 VSUBS 0.00379f
C13516 VDD.n6195 VSUBS 0.0145f
C13517 VDD.t460 VSUBS 0.0114f
C13518 VDD.t462 VSUBS 0.0114f
C13519 VDD.n6196 VSUBS 0.0268f
C13520 VDD.n6197 VSUBS 0.0118f
C13521 VDD.n6198 VSUBS 0.0242f
C13522 VDD.n6199 VSUBS 0.0142f
C13523 VDD.n6200 VSUBS 0.0075f
C13524 VDD.n6201 VSUBS 0.00379f
C13525 VDD.n6202 VSUBS 0.0145f
C13526 VDD.t43 VSUBS 0.0114f
C13527 VDD.t101 VSUBS 0.0114f
C13528 VDD.n6203 VSUBS 0.0268f
C13529 VDD.n6204 VSUBS 0.0118f
C13530 VDD.n6205 VSUBS 0.0242f
C13531 VDD.n6206 VSUBS 0.0142f
C13532 VDD.n6207 VSUBS 0.0075f
C13533 VDD.n6208 VSUBS 0.00379f
C13534 VDD.n6209 VSUBS 0.0202f
C13535 VDD.t7 VSUBS 0.0114f
C13536 VDD.t450 VSUBS 0.0114f
C13537 VDD.n6210 VSUBS 0.0268f
C13538 VDD.n6211 VSUBS 0.0118f
C13539 VDD.n6212 VSUBS 0.0242f
C13540 VDD.n6213 VSUBS 0.0142f
C13541 VDD.n6214 VSUBS 0.215f
C13542 VDD.n6215 VSUBS 0.0867f
C13543 VDD.n6216 VSUBS 0.0867f
C13544 VDD.n6217 VSUBS 0.0867f
C13545 VDD.n6218 VSUBS 0.0867f
C13546 VDD.n6219 VSUBS 0.0867f
C13547 VDD.n6220 VSUBS 0.0867f
C13548 VDD.n6221 VSUBS 0.0867f
C13549 VDD.n6222 VSUBS 0.0867f
C13550 VDD.n6223 VSUBS 0.0867f
C13551 VDD.n6224 VSUBS 0.0867f
C13552 VDD.n6225 VSUBS 0.0867f
C13553 VDD.n6226 VSUBS 0.0867f
C13554 VDD.n6227 VSUBS 0.0867f
C13555 VDD.n6228 VSUBS 0.0867f
C13556 VDD.n6229 VSUBS 0.0867f
C13557 VDD.n6230 VSUBS 0.0867f
C13558 VDD.n6231 VSUBS 0.0867f
C13559 VDD.n6232 VSUBS 0.0867f
C13560 VDD.n6233 VSUBS 0.0867f
C13561 VDD.n6234 VSUBS 0.0867f
C13562 VDD.n6235 VSUBS 0.0867f
C13563 VDD.n6236 VSUBS 0.0867f
C13564 VDD.n6237 VSUBS 0.0867f
C13565 VDD.n6238 VSUBS 0.0867f
C13566 VDD.n6239 VSUBS 0.0867f
C13567 VDD.n6240 VSUBS 0.0867f
C13568 VDD.n6241 VSUBS 0.0867f
C13569 VDD.n6242 VSUBS 0.0867f
C13570 VDD.n6243 VSUBS 0.0867f
C13571 VDD.n6244 VSUBS 0.0867f
C13572 VDD.n6245 VSUBS 0.0867f
C13573 VDD.n6246 VSUBS 0.0867f
C13574 VDD.n6247 VSUBS 0.0867f
C13575 VDD.n6248 VSUBS 0.0867f
C13576 VDD.n6249 VSUBS 0.0867f
C13577 VDD.n6250 VSUBS 0.0867f
C13578 VDD.n6251 VSUBS 0.0867f
C13579 VDD.n6252 VSUBS 0.0867f
C13580 VDD.n6253 VSUBS 0.0198f
C13581 VDD.n6254 VSUBS 0.0277f
C13582 VDD.n6255 VSUBS 0.0198f
C13583 VDD.n6256 VSUBS 0.0448f
C13584 VDD.n6257 VSUBS 0.0155f
C13585 VDD.n6258 VSUBS 0.0217f
C13586 VDD.n6259 VSUBS 0.0408f
C13587 VDD.n6260 VSUBS 0.0198f
C13588 VDD.n6261 VSUBS 0.025f
C13589 VDD.n6262 VSUBS 0.0155f
C13590 VDD.n6263 VSUBS 0.0244f
C13591 VDD.n6264 VSUBS 0.0402f
C13592 VDD.n6265 VSUBS 0.0813f
C13593 VDD.n6266 VSUBS 0.0155f
C13594 VDD.n6267 VSUBS 0.0296f
C13595 VDD.n6268 VSUBS 0.0198f
C13596 VDD.n6269 VSUBS 0.0224f
C13597 VDD.n6270 VSUBS 0.0155f
C13598 VDD.n6271 VSUBS 0.027f
C13599 VDD.n6272 VSUBS 0.0402f
C13600 VDD.n6273 VSUBS 0.0371f
C13601 VDD.n6274 VSUBS 0.0155f
C13602 VDD.n6275 VSUBS 0.0323f
C13603 VDD.n6276 VSUBS 0.0198f
C13604 VDD.n6277 VSUBS 0.0198f
C13605 VDD.n6278 VSUBS 0.0402f
C13606 VDD.n6279 VSUBS 0.0371f
C13607 VDD.n6280 VSUBS 0.0155f
C13608 VDD.n6281 VSUBS 0.0349f
C13609 VDD.n6282 VSUBS 0.0198f
C13610 VDD.n6283 VSUBS 0.0171f
C13611 VDD.n6284 VSUBS 0.0402f
C13612 VDD.n6285 VSUBS 0.0371f
C13613 VDD.n6286 VSUBS 0.0155f
C13614 VDD.n6287 VSUBS 0.0375f
C13615 VDD.n6288 VSUBS 0.0198f
C13616 VDD.n6289 VSUBS 0.0145f
C13617 VDD.n6290 VSUBS 0.0402f
C13618 VDD.n6291 VSUBS 0.0371f
C13619 VDD.n6292 VSUBS 0.0155f
C13620 VDD.n6293 VSUBS 0.0402f
C13621 VDD.n6294 VSUBS 0.0198f
C13622 VDD.n6295 VSUBS 0.0119f
C13623 VDD.n6296 VSUBS 0.0402f
C13624 VDD.n6297 VSUBS 0.0371f
C13625 VDD.n6298 VSUBS 0.0155f
C13626 VDD.n6299 VSUBS 0.0428f
C13627 VDD.n6300 VSUBS 0.0198f
C13628 VDD.n6301 VSUBS 0.00922f
C13629 VDD.n6302 VSUBS 0.0402f
C13630 VDD.n6303 VSUBS 0.0371f
C13631 VDD.n6304 VSUBS 0.0155f
C13632 VDD.n6305 VSUBS 0.0448f
C13633 VDD.n6306 VSUBS 0.0198f
C13634 VDD.n6307 VSUBS 0.00658f
C13635 VDD.n6308 VSUBS 0.0402f
C13636 VDD.n6309 VSUBS 0.0371f
C13637 VDD.n6310 VSUBS 0.0155f
C13638 VDD.n6311 VSUBS 0.0441f
C13639 VDD.n6312 VSUBS 0.0198f
C13640 VDD.n6313 VSUBS 0.0408f
C13641 VDD.n6314 VSUBS 0.00461f
C13642 VDD.n6315 VSUBS 0.0371f
C13643 VDD.n6316 VSUBS 0.0155f
C13644 VDD.n6317 VSUBS 0.0415f
C13645 VDD.n6318 VSUBS 0.0198f
C13646 VDD.n6319 VSUBS 0.0435f
C13647 VDD.n6320 VSUBS 0.00461f
C13648 VDD.n6321 VSUBS 0.0371f
C13649 VDD.n6322 VSUBS 0.0198f
C13650 VDD.n6323 VSUBS 0.0448f
C13651 VDD.n6324 VSUBS 0.0155f
C13652 VDD.n6325 VSUBS 0.00593f
C13653 VDD.n6326 VSUBS 0.0402f
C13654 VDD.n6327 VSUBS 0.0371f
C13655 VDD.n6328 VSUBS 0.0198f
C13656 VDD.n6329 VSUBS 0.0435f
C13657 VDD.n6330 VSUBS 0.0155f
C13658 VDD.n6331 VSUBS 0.00856f
C13659 VDD.n6332 VSUBS 0.0402f
C13660 VDD.n6333 VSUBS 0.0371f
C13661 VDD.n6334 VSUBS 0.0198f
C13662 VDD.n6335 VSUBS 0.0408f
C13663 VDD.n6336 VSUBS 0.0155f
C13664 VDD.n6337 VSUBS 0.0112f
C13665 VDD.n6338 VSUBS 0.0402f
C13666 VDD.n6339 VSUBS 0.0371f
C13667 VDD.n6340 VSUBS 0.0198f
C13668 VDD.n6341 VSUBS 0.0382f
C13669 VDD.n6342 VSUBS 0.0155f
C13670 VDD.n6343 VSUBS 0.0138f
C13671 VDD.n6344 VSUBS 0.0402f
C13672 VDD.n6345 VSUBS 0.0371f
C13673 VDD.n6346 VSUBS 0.0198f
C13674 VDD.n6347 VSUBS 0.0356f
C13675 VDD.n6348 VSUBS 0.0155f
C13676 VDD.n6349 VSUBS 0.0165f
C13677 VDD.n6350 VSUBS 0.0402f
C13678 VDD.n6351 VSUBS 0.0371f
C13679 VDD.n6352 VSUBS 0.0198f
C13680 VDD.n6353 VSUBS 0.0329f
C13681 VDD.n6354 VSUBS 0.0155f
C13682 VDD.n6355 VSUBS 0.0191f
C13683 VDD.n6356 VSUBS 0.0402f
C13684 VDD.n6357 VSUBS 0.0371f
C13685 VDD.n6358 VSUBS 0.0198f
C13686 VDD.n6359 VSUBS 0.0277f
C13687 VDD.n6360 VSUBS 0.0198f
C13688 VDD.n6361 VSUBS 0.0303f
C13689 VDD.n6362 VSUBS 0.0155f
C13690 VDD.n6363 VSUBS 0.0217f
C13691 VDD.n6364 VSUBS 0.0402f
C13692 VDD.n6365 VSUBS 0.0371f
C13693 VDD.n6366 VSUBS 0.0198f
C13694 VDD.n6367 VSUBS 0.025f
C13695 VDD.n6368 VSUBS 0.0155f
C13696 VDD.n6369 VSUBS 0.0244f
C13697 VDD.n6370 VSUBS 0.0402f
C13698 VDD.n6371 VSUBS 0.0371f
C13699 VDD.n6372 VSUBS 0.0155f
C13700 VDD.n6373 VSUBS 0.0296f
C13701 VDD.n6374 VSUBS 0.0198f
C13702 VDD.n6375 VSUBS 0.0224f
C13703 VDD.n6376 VSUBS 0.0155f
C13704 VDD.n6377 VSUBS 0.027f
C13705 VDD.n6378 VSUBS 0.0402f
C13706 VDD.n6379 VSUBS 0.0371f
C13707 VDD.n6380 VSUBS 0.0155f
C13708 VDD.n6381 VSUBS 0.0323f
C13709 VDD.n6382 VSUBS 0.0198f
C13710 VDD.n6383 VSUBS 0.0198f
C13711 VDD.n6384 VSUBS 0.0402f
C13712 VDD.n6385 VSUBS 0.0371f
C13713 VDD.n6386 VSUBS 0.0155f
C13714 VDD.n6387 VSUBS 0.0349f
C13715 VDD.n6388 VSUBS 0.0198f
C13716 VDD.n6389 VSUBS 0.0171f
C13717 VDD.n6390 VSUBS 0.0402f
C13718 VDD.n6391 VSUBS 0.0371f
C13719 VDD.n6392 VSUBS 0.0155f
C13720 VDD.n6393 VSUBS 0.0375f
C13721 VDD.n6394 VSUBS 0.0198f
C13722 VDD.n6395 VSUBS 0.0145f
C13723 VDD.n6396 VSUBS 0.0402f
C13724 VDD.n6397 VSUBS 0.0371f
C13725 VDD.n6398 VSUBS 0.0155f
C13726 VDD.n6399 VSUBS 0.0402f
C13727 VDD.n6400 VSUBS 0.0198f
C13728 VDD.n6401 VSUBS 0.0119f
C13729 VDD.n6402 VSUBS 0.0402f
C13730 VDD.n6403 VSUBS 0.0371f
C13731 VDD.n6404 VSUBS 0.0155f
C13732 VDD.n6405 VSUBS 0.0428f
C13733 VDD.n6406 VSUBS 0.0198f
C13734 VDD.n6407 VSUBS 0.00922f
C13735 VDD.n6408 VSUBS 0.0402f
C13736 VDD.n6409 VSUBS 0.0371f
C13737 VDD.n6410 VSUBS 0.0155f
C13738 VDD.n6411 VSUBS 0.0448f
C13739 VDD.n6412 VSUBS 0.0198f
C13740 VDD.n6413 VSUBS 0.00658f
C13741 VDD.n6414 VSUBS 0.0402f
C13742 VDD.n6415 VSUBS 0.0371f
C13743 VDD.n6416 VSUBS 0.0155f
C13744 VDD.n6417 VSUBS 0.0441f
C13745 VDD.n6418 VSUBS 0.0198f
C13746 VDD.n6419 VSUBS 0.0408f
C13747 VDD.n6420 VSUBS 0.00461f
C13748 VDD.n6421 VSUBS 0.0371f
C13749 VDD.n6422 VSUBS 0.0327f
C13750 VDD.n6423 VSUBS 0.0415f
C13751 VDD.n6424 VSUBS 0.0198f
C13752 VDD.n6425 VSUBS 0.0435f
C13753 VDD.n6426 VSUBS 0.00461f
C13754 VDD.n6427 VSUBS 0.0371f
C13755 VDD.n6428 VSUBS 0.0198f
C13756 VDD.n6429 VSUBS 0.0461f
C13757 VDD.n6430 VSUBS 0.0448f
C13758 VDD.n6431 VSUBS 0.0371f
C13759 VDD.n6432 VSUBS 0.0421f
C13760 VDD.n6433 VSUBS 0.0421f
C13761 VDD.n6434 VSUBS 0.0421f
C13762 VDD.n6435 VSUBS 0.0421f
C13763 VDD.n6436 VSUBS 0.0421f
C13764 VDD.n6437 VSUBS 0.0421f
C13765 VDD.n6438 VSUBS 0.0421f
C13766 VDD.n6439 VSUBS 0.0421f
C13767 VDD.n6440 VSUBS 0.0421f
C13768 VDD.n6441 VSUBS 0.0421f
C13769 VDD.n6442 VSUBS 0.0421f
C13770 VDD.n6443 VSUBS 0.0421f
C13771 VDD.n6444 VSUBS 0.0421f
C13772 VDD.n6445 VSUBS 0.0421f
C13773 VDD.n6446 VSUBS 0.0421f
C13774 VDD.n6447 VSUBS 0.0421f
C13775 VDD.n6448 VSUBS 0.0421f
C13776 VDD.n6449 VSUBS 0.0421f
C13777 VDD.n6450 VSUBS 0.0421f
C13778 VDD.n6451 VSUBS 0.0421f
C13779 VDD.n6452 VSUBS 0.0421f
C13780 VDD.n6453 VSUBS 0.0421f
C13781 VDD.n6454 VSUBS 0.0421f
C13782 VDD.n6455 VSUBS 0.0421f
C13783 VDD.n6456 VSUBS 0.0421f
C13784 VDD.n6457 VSUBS 0.0421f
C13785 VDD.n6458 VSUBS 0.0421f
C13786 VDD.n6459 VSUBS 0.0421f
C13787 VDD.n6460 VSUBS 0.0421f
C13788 VDD.n6461 VSUBS 0.0421f
C13789 VDD.n6462 VSUBS 0.0421f
C13790 VDD.n6463 VSUBS 0.0421f
C13791 VDD.n6464 VSUBS 0.0421f
C13792 VDD.n6465 VSUBS 0.0198f
C13793 VDD.n6466 VSUBS 0.0421f
C13794 VDD.n6467 VSUBS 0.0421f
C13795 VDD.n6468 VSUBS 0.0198f
C13796 VDD.n6469 VSUBS 0.0421f
C13797 VDD.n6470 VSUBS 0.0155f
C13798 VDD.n6471 VSUBS 0.0421f
C13799 VDD.n6472 VSUBS 0.0198f
C13800 VDD.n6473 VSUBS 0.0421f
C13801 VDD.n6474 VSUBS 0.0155f
C13802 VDD.n6475 VSUBS 0.0421f
C13803 VDD.n6476 VSUBS 0.0198f
C13804 VDD.n6477 VSUBS 0.0421f
C13805 VDD.n6478 VSUBS 0.0155f
C13806 VDD.n6479 VSUBS 0.0421f
C13807 VDD.n6480 VSUBS 0.0198f
C13808 VDD.n6481 VSUBS 0.0421f
C13809 VDD.n6482 VSUBS 0.0325f
C13810 VDD.n6483 VSUBS 0.0421f
C13811 VDD.n6484 VSUBS 0.0198f
C13812 VDD.n6485 VSUBS 0.0502f
C13813 VDD.n6486 VSUBS 0.0198f
C13814 VDD.n6487 VSUBS 0.0198f
C13815 VDD.n6489 VSUBS 0.0198f
C13816 VDD.n6490 VSUBS 0.0287f
C13817 VDD.n6492 VSUBS 0.0672f
C13818 VDD.n6494 VSUBS 0.0333f
C13819 VDD.n6495 VSUBS 0.0896f
C13820 VDD.n6496 VSUBS 0.0198f
C13821 VDD.n6497 VSUBS 0.0481f
C13822 VDD.n6498 VSUBS 0.064f
C13823 VDD.n6500 VSUBS 0.0198f
C13824 VDD.n6501 VSUBS 0.0777f
C13825 VDD.n6502 VSUBS 0.0198f
C13826 VDD.n6503 VSUBS 0.0474f
C13827 VDD.n6504 VSUBS 0.0448f
C13828 VDD.n6505 VSUBS 1.51f
C13829 VDD.n6506 VSUBS 0.0421f
C13830 VDD.n6507 VSUBS 0.0421f
C13831 VDD.n6508 VSUBS 0.0421f
C13832 VDD.n6509 VSUBS 0.0421f
C13833 VDD.n6510 VSUBS 0.0421f
C13834 VDD.n6511 VSUBS 0.0421f
C13835 VDD.n6512 VSUBS 0.0421f
C13836 VDD.n6513 VSUBS 0.0421f
C13837 VDD.n6514 VSUBS 0.0421f
C13838 VDD.n6515 VSUBS 0.0421f
C13839 VDD.n6516 VSUBS 0.0421f
C13840 VDD.n6517 VSUBS 0.0421f
C13841 VDD.n6518 VSUBS 0.0421f
C13842 VDD.n6519 VSUBS 0.0421f
C13843 VDD.n6520 VSUBS 0.0421f
C13844 VDD.n6521 VSUBS 0.0421f
C13845 VDD.n6522 VSUBS 0.0421f
C13846 VDD.n6523 VSUBS 0.0421f
C13847 VDD.n6524 VSUBS 0.0421f
C13848 VDD.n6525 VSUBS 0.0421f
C13849 VDD.n6526 VSUBS 0.0421f
C13850 VDD.n6527 VSUBS 0.0421f
C13851 VDD.n6528 VSUBS 0.0421f
C13852 VDD.n6529 VSUBS 0.0421f
C13853 VDD.n6530 VSUBS 0.0421f
C13854 VDD.n6531 VSUBS 0.0421f
C13855 VDD.n6532 VSUBS 0.0421f
C13856 VDD.n6533 VSUBS 0.0421f
C13857 VDD.n6534 VSUBS 0.0421f
C13858 VDD.n6535 VSUBS 0.0421f
C13859 VDD.n6536 VSUBS 0.0421f
C13860 VDD.n6537 VSUBS 0.0421f
C13861 VDD.n6538 VSUBS 0.0421f
C13862 VDD.n6539 VSUBS 0.0421f
C13863 VDD.n6540 VSUBS 0.0421f
C13864 VDD.n6541 VSUBS 0.0421f
C13865 VDD.n6542 VSUBS 0.0421f
C13866 VDD.n6543 VSUBS 0.0421f
C13867 VDD.n6544 VSUBS 0.0421f
C13868 VDD.n6545 VSUBS 0.0421f
C13869 VDD.n6546 VSUBS 0.0421f
C13870 VDD.n6547 VSUBS 0.0421f
C13871 VDD.n6548 VSUBS 0.0421f
C13872 VDD.n6549 VSUBS 0.0421f
C13873 VDD.n6550 VSUBS 0.0421f
C13874 VDD.n6551 VSUBS 0.0421f
C13875 VDD.n6552 VSUBS 0.0421f
C13876 VDD.n6553 VSUBS 0.0421f
C13877 VDD.n6554 VSUBS 0.0421f
C13878 VDD.n6555 VSUBS 0.0421f
C13879 VDD.n6556 VSUBS 0.0421f
C13880 VDD.n6557 VSUBS 0.0421f
C13881 VDD.n6558 VSUBS 0.0421f
C13882 VDD.n6559 VSUBS 0.0421f
C13883 VDD.n6560 VSUBS 0.0421f
C13884 VDD.n6561 VSUBS 0.0421f
C13885 VDD.n6562 VSUBS 0.0421f
C13886 VDD.n6563 VSUBS 0.0421f
C13887 VDD.n6564 VSUBS 0.0421f
C13888 VDD.n6565 VSUBS 0.0421f
C13889 VDD.n6566 VSUBS 0.0421f
C13890 VDD.n6567 VSUBS 0.0421f
C13891 VDD.n6568 VSUBS 0.0421f
C13892 VDD.n6569 VSUBS 0.0421f
C13893 VDD.n6570 VSUBS 0.0421f
C13894 VDD.n6571 VSUBS 0.0421f
C13895 VDD.n6572 VSUBS 0.0421f
C13896 VDD.n6573 VSUBS 0.0198f
C13897 VDD.n6574 VSUBS 0.0421f
C13898 VDD.n6575 VSUBS 0.0421f
C13899 VDD.n6576 VSUBS 0.0198f
C13900 VDD.n6577 VSUBS 0.0421f
C13901 VDD.n6578 VSUBS 0.0155f
C13902 VDD.n6579 VSUBS 0.0421f
C13903 VDD.n6580 VSUBS 0.0198f
C13904 VDD.n6581 VSUBS 0.0421f
C13905 VDD.n6582 VSUBS 0.0155f
C13906 VDD.n6583 VSUBS 0.0421f
C13907 VDD.n6584 VSUBS 0.0198f
C13908 VDD.n6585 VSUBS 0.0421f
C13909 VDD.n6586 VSUBS 0.0155f
C13910 VDD.n6587 VSUBS 0.0421f
C13911 VDD.n6588 VSUBS 0.0198f
C13912 VDD.n6589 VSUBS 0.0421f
C13913 VDD.n6590 VSUBS 0.0155f
C13914 VDD.n6591 VSUBS 0.0421f
C13915 VDD.n6592 VSUBS 0.0198f
C13916 VDD.n6593 VSUBS 0.0421f
C13917 VDD.n6594 VSUBS 0.0155f
C13918 VDD.n6595 VSUBS 0.0421f
C13919 VDD.n6596 VSUBS 0.0198f
C13920 VDD.n6597 VSUBS 0.0421f
C13921 VDD.n6598 VSUBS 0.0155f
C13922 VDD.n6599 VSUBS 0.0421f
C13923 VDD.n6600 VSUBS 0.0198f
C13924 VDD.n6601 VSUBS 0.0421f
C13925 VDD.n6602 VSUBS 0.0155f
C13926 VDD.n6603 VSUBS 0.0421f
C13927 VDD.n6604 VSUBS 0.0198f
C13928 VDD.n6605 VSUBS 0.0421f
C13929 VDD.n6606 VSUBS 0.0155f
C13930 VDD.n6607 VSUBS 0.0421f
C13931 VDD.n6608 VSUBS 0.0198f
C13932 VDD.n6609 VSUBS 0.0421f
C13933 VDD.n6610 VSUBS 0.0155f
C13934 VDD.n6611 VSUBS 0.0421f
C13935 VDD.n6612 VSUBS 0.0198f
C13936 VDD.n6613 VSUBS 0.0421f
C13937 VDD.n6614 VSUBS 0.0155f
C13938 VDD.n6615 VSUBS 0.0421f
C13939 VDD.n6616 VSUBS 0.0198f
C13940 VDD.n6617 VSUBS 0.0421f
C13941 VDD.n6618 VSUBS 0.0155f
C13942 VDD.n6619 VSUBS 0.0421f
C13943 VDD.n6620 VSUBS 0.0198f
C13944 VDD.n6621 VSUBS 0.039f
C13945 VDD.n6622 VSUBS 0.0421f
C13946 VDD.n6623 VSUBS 0.0421f
C13947 VDD.n6624 VSUBS 0.0421f
C13948 VDD.n6625 VSUBS 0.0421f
C13949 VDD.n6626 VSUBS 0.0421f
C13950 VDD.n6627 VSUBS 0.0421f
C13951 VDD.n6628 VSUBS 0.0421f
C13952 VDD.n6629 VSUBS 0.0421f
C13953 VDD.n6630 VSUBS 0.0421f
C13954 VDD.n6631 VSUBS 0.0421f
C13955 VDD.n6632 VSUBS 0.0421f
C13956 VDD.n6633 VSUBS 0.0421f
C13957 VDD.n6634 VSUBS 0.0421f
C13958 VDD.n6635 VSUBS 0.0421f
C13959 VDD.n6636 VSUBS 0.0421f
C13960 VDD.n6637 VSUBS 0.0421f
C13961 VDD.n6638 VSUBS 0.0421f
C13962 VDD.n6639 VSUBS 0.0421f
C13963 VDD.n6640 VSUBS 0.0421f
C13964 VDD.n6641 VSUBS 0.0421f
C13965 VDD.n6642 VSUBS 0.0421f
C13966 VDD.n6643 VSUBS 0.0421f
C13967 VDD.n6644 VSUBS 0.0421f
C13968 VDD.n6645 VSUBS 0.0421f
C13969 VDD.n6646 VSUBS 0.0421f
C13970 VDD.n6647 VSUBS 0.0421f
C13971 VDD.n6648 VSUBS 0.0421f
C13972 VDD.n6649 VSUBS 0.0421f
C13973 VDD.n6650 VSUBS 0.0421f
C13974 VDD.n6651 VSUBS 0.0421f
C13975 VDD.n6652 VSUBS 0.0198f
C13976 VDD.n6653 VSUBS 0.0421f
C13977 VDD.n6654 VSUBS 0.0155f
C13978 VDD.n6655 VSUBS 0.0421f
C13979 VDD.n6656 VSUBS 0.0198f
C13980 VDD.n6657 VSUBS 0.0421f
C13981 VDD.n6658 VSUBS 0.0155f
C13982 VDD.n6659 VSUBS 0.0421f
C13983 VDD.n6660 VSUBS 0.0198f
C13984 VDD.n6661 VSUBS 0.0421f
C13985 VDD.n6662 VSUBS 0.0155f
C13986 VDD.n6663 VSUBS 0.0421f
C13987 VDD.n6664 VSUBS 0.0198f
C13988 VDD.n6665 VSUBS 0.0421f
C13989 VDD.n6666 VSUBS 0.0155f
C13990 VDD.n6667 VSUBS 0.0421f
C13991 VDD.n6668 VSUBS 0.0198f
C13992 VDD.n6669 VSUBS 0.0421f
C13993 VDD.n6670 VSUBS 0.0155f
C13994 VDD.n6671 VSUBS 0.0421f
C13995 VDD.n6672 VSUBS 0.0198f
C13996 VDD.n6673 VSUBS 0.0421f
C13997 VDD.n6674 VSUBS 0.0155f
C13998 VDD.n6675 VSUBS 0.0421f
C13999 VDD.n6676 VSUBS 0.0198f
C14000 VDD.n6677 VSUBS 0.0421f
C14001 VDD.n6678 VSUBS 0.0155f
C14002 VDD.n6679 VSUBS 0.0421f
C14003 VDD.n6680 VSUBS 0.0198f
C14004 VDD.n6681 VSUBS 0.0421f
C14005 VDD.n6682 VSUBS 0.0155f
C14006 VDD.n6683 VSUBS 0.0421f
C14007 VDD.n6684 VSUBS 0.0198f
C14008 VDD.n6685 VSUBS 0.0421f
C14009 VDD.n6686 VSUBS 0.0155f
C14010 VDD.n6687 VSUBS 0.0421f
C14011 VDD.n6688 VSUBS 0.0198f
C14012 VDD.n6689 VSUBS 0.0421f
C14013 VDD.n6690 VSUBS 0.0155f
C14014 VDD.n6691 VSUBS 0.0421f
C14015 VDD.n6692 VSUBS 0.0198f
C14016 VDD.n6693 VSUBS 0.0421f
C14017 VDD.n6694 VSUBS 0.0155f
C14018 VDD.n6695 VSUBS 0.0341f
C14019 VDD.n6696 VSUBS 9.03f
C14020 VDD.n6697 VSUBS 0.401f
C14021 VDD.n6698 VSUBS 1.89f
C14022 VDD.n6699 VSUBS 0.457f
C14023 VDD.n6700 VSUBS 0.454f
C14024 VDD.n6701 VSUBS 0.447f
C14025 VDD.n6702 VSUBS 0.349f
C14026 VDD.n6703 VSUBS 0.276f
C14027 VDD.n6704 VSUBS 0.441f
C14028 VDD.n6705 VSUBS 0.452f
C14029 VDD.n6706 VSUBS 0.452f
C14030 VDD.n6707 VSUBS 0.452f
C14031 VDD.n6708 VSUBS 0.458f
C14032 VDD.n6709 VSUBS 0.318f
C14033 VDD.n6710 VSUBS 0.0466f
C14034 VDD.n6711 VSUBS 0.0842f
C14035 VDD.n6712 VSUBS 0.0198f
C14036 VDD.n6713 VSUBS 0.052f
C14037 VDD.n6714 VSUBS 0.0842f
C14038 VDD.n6715 VSUBS 0.0198f
C14039 VDD.n6716 VSUBS 0.0738f
C14040 VDD.n6717 VSUBS 0.0842f
C14041 VDD.n6718 VSUBS 0.0198f
C14042 VDD.n6719 VSUBS 0.0441f
C14043 VDD.n6720 VSUBS 0.0842f
C14044 VDD.n6721 VSUBS 0.0198f
C14045 VDD.n6722 VSUBS 0.0441f
C14046 VDD.n6723 VSUBS 0.0842f
C14047 VDD.n6724 VSUBS 0.0198f
C14048 VDD.n6725 VSUBS 0.0441f
C14049 VDD.n6726 VSUBS 0.0842f
C14050 VDD.n6727 VSUBS 0.0198f
C14051 VDD.n6728 VSUBS 0.0441f
C14052 VDD.n6729 VSUBS 0.0842f
C14053 VDD.n6730 VSUBS 0.0198f
C14054 VDD.n6731 VSUBS 0.0441f
C14055 VDD.n6732 VSUBS 0.0842f
C14056 VDD.n6733 VSUBS 0.0198f
C14057 VDD.n6734 VSUBS 0.0441f
C14058 VDD.n6735 VSUBS 0.0842f
C14059 VDD.n6736 VSUBS 0.0198f
C14060 VDD.n6737 VSUBS 0.0441f
C14061 VDD.n6738 VSUBS 0.0842f
C14062 VDD.n6739 VSUBS 0.0198f
C14063 VDD.n6740 VSUBS 0.0441f
C14064 VDD.n6741 VSUBS 0.0842f
C14065 VDD.n6742 VSUBS 0.0198f
C14066 VDD.n6743 VSUBS 0.0441f
C14067 VDD.n6744 VSUBS 0.0842f
C14068 VDD.n6745 VSUBS 0.0198f
C14069 VDD.n6746 VSUBS 0.0441f
C14070 VDD.n6747 VSUBS 0.0842f
C14071 VDD.n6748 VSUBS 0.0198f
C14072 VDD.n6749 VSUBS 0.0499f
C14073 VDD.n6750 VSUBS 0.0842f
C14074 VDD.n6751 VSUBS 0.0198f
C14075 VDD.n6752 VSUBS 0.0899f
C14076 VDD.n6753 VSUBS 0.0842f
C14077 VDD.n6754 VSUBS 0.0198f
C14078 VDD.n6755 VSUBS 0.0858f
C14079 VDD.n6756 VSUBS 0.0842f
C14080 VDD.n6757 VSUBS 0.0198f
C14081 VDD.n6758 VSUBS 0.0858f
C14082 VDD.n6759 VSUBS 0.0842f
C14083 VDD.n6760 VSUBS 0.0198f
C14084 VDD.n6761 VSUBS 0.0858f
C14085 VDD.n6762 VSUBS 0.0842f
C14086 VDD.n6763 VSUBS 0.0198f
C14087 VDD.n6764 VSUBS 0.0858f
C14088 VDD.n6765 VSUBS 0.0842f
C14089 VDD.n6766 VSUBS 0.0198f
C14090 VDD.n6767 VSUBS 0.0858f
C14091 VDD.n6768 VSUBS 0.0842f
C14092 VDD.n6769 VSUBS 0.0198f
C14093 VDD.n6770 VSUBS 0.0858f
C14094 VDD.n6771 VSUBS 0.0842f
C14095 VDD.n6772 VSUBS 0.0198f
C14096 VDD.n6773 VSUBS 0.0858f
C14097 VDD.n6774 VSUBS 0.0842f
C14098 VDD.n6775 VSUBS 0.0198f
C14099 VDD.n6776 VSUBS 0.0858f
C14100 VDD.n6777 VSUBS 0.0842f
C14101 VDD.n6778 VSUBS 0.0198f
C14102 VDD.n6779 VSUBS 0.0858f
C14103 VDD.n6780 VSUBS 0.0842f
C14104 VDD.n6781 VSUBS 0.0198f
C14105 VDD.n6782 VSUBS 0.0656f
C14106 VDD.n6783 VSUBS 0.0434f
C14107 VDD.n6784 VSUBS 0.0842f
C14108 VDD.n6785 VSUBS 0.0198f
C14109 VDD.n6786 VSUBS 0.0647f
C14110 VDD.n6787 VSUBS 0.0842f
C14111 VDD.n6788 VSUBS 0.0198f
C14112 VDD.n6789 VSUBS 0.0607f
C14113 VDD.n6790 VSUBS 0.0448f
C14114 VDD.n6791 VSUBS 0.644f
C14115 pdrv1.n0 VSUBS 4.46f
C14116 pdrv1.n1 VSUBS 1.27f
C14117 pdrv1.n2 VSUBS 1.27f
C14118 pdrv1.n3 VSUBS 1.27f
C14119 pdrv1.n4 VSUBS 1.27f
C14120 pdrv1.n5 VSUBS 1.27f
C14121 pdrv1.n6 VSUBS 1.27f
C14122 pdrv1.n7 VSUBS 1.27f
C14123 pdrv1.n8 VSUBS 1.27f
C14124 pdrv1.n9 VSUBS 1.29f
C14125 pdrv1.n10 VSUBS 1.32f
C14126 pdrv1.n11 VSUBS 1.29f
C14127 pdrv1.n12 VSUBS 1.29f
C14128 pdrv1.n13 VSUBS 1.29f
C14129 pdrv1.n14 VSUBS 1.29f
C14130 pdrv1.n15 VSUBS 1.29f
C14131 pdrv1.n16 VSUBS 1.29f
C14132 pdrv1.n17 VSUBS 1.29f
C14133 pdrv1.n18 VSUBS 1.29f
C14134 pdrv1.n19 VSUBS 1.32f
C14135 pdrv1.n20 VSUBS 1.31f
C14136 pdrv1.n21 VSUBS 1.28f
C14137 pdrv1.n22 VSUBS 1.28f
C14138 pdrv1.n23 VSUBS 1.28f
C14139 pdrv1.n24 VSUBS 1.28f
C14140 pdrv1.n25 VSUBS 1.28f
C14141 pdrv1.n26 VSUBS 1.28f
C14142 pdrv1.n27 VSUBS 1.28f
C14143 pdrv1.n28 VSUBS 1.28f
C14144 pdrv1.n29 VSUBS 4.86f
C14145 pdrv1.n30 VSUBS 2.62f
C14146 pdrv1.n31 VSUBS 0.339f
C14147 pdrv1.n32 VSUBS 0.339f
C14148 pdrv1.n33 VSUBS 0.351f
C14149 pdrv1.n34 VSUBS 0.657f
C14150 pdrv1.n35 VSUBS 0.675f
C14151 pdrv1.n36 VSUBS 0.657f
C14152 pdrv1.n37 VSUBS 0.657f
C14153 pdrv1.n38 VSUBS 0.657f
C14154 pdrv1.n39 VSUBS 0.657f
C14155 pdrv1.n40 VSUBS 0.657f
C14156 pdrv1.n41 VSUBS 0.657f
C14157 pdrv1.n42 VSUBS 0.657f
C14158 pdrv1.n43 VSUBS 0.657f
C14159 pdrv1.n44 VSUBS 0.657f
C14160 pdrv1.n45 VSUBS 0.657f
C14161 pdrv1.n46 VSUBS 0.657f
C14162 pdrv1.n47 VSUBS 0.657f
C14163 pdrv1.n48 VSUBS 0.657f
C14164 pdrv1.n49 VSUBS 0.657f
C14165 pdrv1.n50 VSUBS 0.657f
C14166 pdrv1.n51 VSUBS 0.657f
C14167 pdrv1.n52 VSUBS 0.657f
C14168 pdrv1.n53 VSUBS 0.675f
C14169 pdrv1.t141 VSUBS 0.142f
C14170 pdrv1.t43 VSUBS 0.142f
C14171 pdrv1.t132 VSUBS 0.142f
C14172 pdrv1.t33 VSUBS 0.142f
C14173 pdrv1.t44 VSUBS 0.142f
C14174 pdrv1.t194 VSUBS 0.142f
C14175 pdrv1.t112 VSUBS 0.142f
C14176 pdrv1.t61 VSUBS 0.142f
C14177 pdrv1.t163 VSUBS 0.142f
C14178 pdrv1.t173 VSUBS 0.142f
C14179 pdrv1.t90 VSUBS 0.142f
C14180 pdrv1.t35 VSUBS 0.142f
C14181 pdrv1.t186 VSUBS 0.142f
C14182 pdrv1.t107 VSUBS 0.142f
C14183 pdrv1.t41 VSUBS 0.142f
C14184 pdrv1.t168 VSUBS 0.142f
C14185 pdrv1.t12 VSUBS 0.142f
C14186 pdrv1.t63 VSUBS 0.142f
C14187 pdrv1.t154 VSUBS 0.142f
C14188 pdrv1.t146 VSUBS 0.142f
C14189 pdrv1.t45 VSUBS 0.142f
C14190 pdrv1.t108 VSUBS 0.142f
C14191 pdrv1.t188 VSUBS 0.142f
C14192 pdrv1.t36 VSUBS 0.142f
C14193 pdrv1.t30 VSUBS 0.142f
C14194 pdrv1.t130 VSUBS 0.142f
C14195 pdrv1.t166 VSUBS 0.142f
C14196 pdrv1.t135 VSUBS 0.142f
C14197 pdrv1.t174 VSUBS 0.142f
C14198 pdrv1.t16 VSUBS 0.142f
C14199 pdrv1.t66 VSUBS 0.142f
C14200 pdrv1.t115 VSUBS 0.142f
C14201 pdrv1.t200 VSUBS 0.142f
C14202 pdrv1.t125 VSUBS 0.142f
C14203 pdrv1.t156 VSUBS 0.142f
C14204 pdrv1.t199 VSUBS 0.142f
C14205 pdrv1.t50 VSUBS 0.142f
C14206 pdrv1.t144 VSUBS 0.142f
C14207 pdrv1.t182 VSUBS 0.142f
C14208 pdrv1.t27 VSUBS 0.142f
C14209 pdrv1.t5 VSUBS 0.142f
C14210 pdrv1.t121 VSUBS 0.142f
C14211 pdrv1.t196 VSUBS 0.142f
C14212 pdrv1.t113 VSUBS 0.142f
C14213 pdrv1.t122 VSUBS 0.142f
C14214 pdrv1.t76 VSUBS 0.142f
C14215 pdrv1.t171 VSUBS 0.142f
C14216 pdrv1.t133 VSUBS 0.142f
C14217 pdrv1.t39 VSUBS 0.142f
C14218 pdrv1.t51 VSUBS 0.142f
C14219 pdrv1.t151 VSUBS 0.142f
C14220 pdrv1.t116 VSUBS 0.142f
C14221 pdrv1.t67 VSUBS 0.142f
C14222 pdrv1.t165 VSUBS 0.142f
C14223 pdrv1.t120 VSUBS 0.142f
C14224 pdrv1.t46 VSUBS 0.142f
C14225 pdrv1.t95 VSUBS 0.142f
C14226 pdrv1.t134 VSUBS 0.142f
C14227 pdrv1.t22 VSUBS 0.142f
C14228 pdrv1.t15 VSUBS 0.142f
C14229 pdrv1.t123 VSUBS 0.142f
C14230 pdrv1.t167 VSUBS 0.142f
C14231 pdrv1.t68 VSUBS 0.142f
C14232 pdrv1.t117 VSUBS 0.142f
C14233 pdrv1.t111 VSUBS 0.142f
C14234 pdrv1.t192 VSUBS 0.142f
C14235 pdrv1.t40 VSUBS 0.142f
C14236 pdrv1.t201 VSUBS 0.142f
C14237 pdrv1.t52 VSUBS 0.142f
C14238 pdrv1.t99 VSUBS 0.142f
C14239 pdrv1.t138 VSUBS 0.142f
C14240 pdrv1.t176 VSUBS 0.142f
C14241 pdrv1.t82 VSUBS 0.142f
C14242 pdrv1.t183 VSUBS 0.142f
C14243 pdrv1.t28 VSUBS 0.142f
C14244 pdrv1.t80 VSUBS 0.142f
C14245 pdrv1.t126 VSUBS 0.142f
C14246 pdrv1.t9 VSUBS 0.142f
C14247 pdrv1.t60 VSUBS 0.142f
C14248 pdrv1.t109 VSUBS 0.142f
C14249 pdrv1.n54 VSUBS 2.52f
C14250 pdrv1.t158 VSUBS 0.142f
C14251 pdrv1.t72 VSUBS 0.142f
C14252 pdrv1.t153 VSUBS 0.142f
C14253 pdrv1.t62 VSUBS 0.142f
C14254 pdrv1.t74 VSUBS 0.142f
C14255 pdrv1.t20 VSUBS 0.142f
C14256 pdrv1.t131 VSUBS 0.142f
C14257 pdrv1.t91 VSUBS 0.142f
C14258 pdrv1.t189 VSUBS 0.142f
C14259 pdrv1.t197 VSUBS 0.142f
C14260 pdrv1.t114 VSUBS 0.142f
C14261 pdrv1.t64 VSUBS 0.142f
C14262 pdrv1.t13 VSUBS 0.142f
C14263 pdrv1.t128 VSUBS 0.142f
C14264 pdrv1.t71 VSUBS 0.142f
C14265 pdrv1.t193 VSUBS 0.142f
C14266 pdrv1.t42 VSUBS 0.142f
C14267 pdrv1.t94 VSUBS 0.142f
C14268 pdrv1.t106 VSUBS 0.142f
C14269 pdrv1.t178 VSUBS 0.142f
C14270 pdrv1.t185 VSUBS 0.142f
C14271 pdrv1.t169 VSUBS 0.142f
C14272 pdrv1.t181 VSUBS 0.142f
C14273 pdrv1.t75 VSUBS 0.142f
C14274 pdrv1.t88 VSUBS 0.142f
C14275 pdrv1.t129 VSUBS 0.142f
C14276 pdrv1.t140 VSUBS 0.142f
C14277 pdrv1.t14 VSUBS 0.142f
C14278 pdrv1.t31 VSUBS 0.142f
C14279 pdrv1.t65 VSUBS 0.142f
C14280 pdrv1.t83 VSUBS 0.142f
C14281 pdrv1.t58 VSUBS 0.142f
C14282 pdrv1.t73 VSUBS 0.142f
C14283 pdrv1.t149 VSUBS 0.142f
C14284 pdrv1.t159 VSUBS 0.142f
C14285 pdrv1.t190 VSUBS 0.142f
C14286 pdrv1.t4 VSUBS 0.142f
C14287 pdrv1.t155 VSUBS 0.142f
C14288 pdrv1.t164 VSUBS 0.142f
C14289 pdrv1.t198 VSUBS 0.142f
C14290 pdrv1.t11 VSUBS 0.142f
C14291 pdrv1.t49 VSUBS 0.142f
C14292 pdrv1.t59 VSUBS 0.142f
C14293 pdrv1.t98 VSUBS 0.142f
C14294 pdrv1.t110 VSUBS 0.142f
C14295 pdrv1.t137 VSUBS 0.142f
C14296 pdrv1.t145 VSUBS 0.142f
C14297 pdrv1.t26 VSUBS 0.142f
C14298 pdrv1.t38 VSUBS 0.142f
C14299 pdrv1.t143 VSUBS 0.142f
C14300 pdrv1.t150 VSUBS 0.142f
C14301 pdrv1.t180 VSUBS 0.142f
C14302 pdrv1.t191 VSUBS 0.142f
C14303 pdrv1.t25 VSUBS 0.142f
C14304 pdrv1.t37 VSUBS 0.142f
C14305 pdrv1.t79 VSUBS 0.142f
C14306 pdrv1.t92 VSUBS 0.142f
C14307 pdrv1.t162 VSUBS 0.142f
C14308 pdrv1.t175 VSUBS 0.142f
C14309 pdrv1.t8 VSUBS 0.142f
C14310 pdrv1.t21 VSUBS 0.142f
C14311 pdrv1.t57 VSUBS 0.142f
C14312 pdrv1.t70 VSUBS 0.142f
C14313 pdrv1.n55 VSUBS 0.256f
C14314 pdrv1.t118 VSUBS 0.142f
C14315 pdrv1.t17 VSUBS 0.142f
C14316 pdrv1.t23 VSUBS 0.142f
C14317 pdrv1.t136 VSUBS 0.142f
C14318 pdrv1.t96 VSUBS 0.142f
C14319 pdrv1.t47 VSUBS 0.142f
C14320 pdrv1.t147 VSUBS 0.142f
C14321 pdrv1.t100 VSUBS 0.142f
C14322 pdrv1.t19 VSUBS 0.142f
C14323 pdrv1.t69 VSUBS 0.142f
C14324 pdrv1.t119 VSUBS 0.142f
C14325 pdrv1.t2 VSUBS 0.142f
C14326 pdrv1.t195 VSUBS 0.142f
C14327 pdrv1.t103 VSUBS 0.142f
C14328 pdrv1.t148 VSUBS 0.142f
C14329 pdrv1.t48 VSUBS 0.142f
C14330 pdrv1.t97 VSUBS 0.142f
C14331 pdrv1.t89 VSUBS 0.142f
C14332 pdrv1.t172 VSUBS 0.142f
C14333 pdrv1.t18 VSUBS 0.142f
C14334 pdrv1.t179 VSUBS 0.142f
C14335 pdrv1.t24 VSUBS 0.142f
C14336 pdrv1.t77 VSUBS 0.142f
C14337 pdrv1.t124 VSUBS 0.142f
C14338 pdrv1.t157 VSUBS 0.142f
C14339 pdrv1.t56 VSUBS 0.142f
C14340 pdrv1.t160 VSUBS 0.142f
C14341 pdrv1.t6 VSUBS 0.142f
C14342 pdrv1.t54 VSUBS 0.142f
C14343 pdrv1.t105 VSUBS 0.142f
C14344 pdrv1.t187 VSUBS 0.142f
C14345 pdrv1.t34 VSUBS 0.142f
C14346 pdrv1.t87 VSUBS 0.142f
C14347 pdrv1.t55 VSUBS 0.142f
C14348 pdrv1.t7 VSUBS 0.142f
C14349 pdrv1.t84 VSUBS 0.142f
C14350 pdrv1.t139 VSUBS 0.142f
C14351 pdrv1.t29 VSUBS 0.142f
C14352 pdrv1.t81 VSUBS 0.142f
C14353 pdrv1.t127 VSUBS 0.142f
C14354 pdrv1.t10 VSUBS 0.142f
C14355 pdrv1.t3 VSUBS 0.142f
C14356 pdrv1.t104 VSUBS 0.142f
C14357 pdrv1.t142 VSUBS 0.142f
C14358 pdrv1.t32 VSUBS 0.142f
C14359 pdrv1.t86 VSUBS 0.142f
C14360 pdrv1.t78 VSUBS 0.142f
C14361 pdrv1.t161 VSUBS 0.142f
C14362 pdrv1.t85 VSUBS 0.142f
C14363 pdrv1.t170 VSUBS 0.142f
C14364 pdrv1.n56 VSUBS 0.238f
C14365 pdrv1.t184 VSUBS 0.142f
C14366 pdrv1.t101 VSUBS 0.142f
C14367 pdrv1.t177 VSUBS 0.142f
C14368 pdrv1.t93 VSUBS 0.142f
C14369 pdrv1.t102 VSUBS 0.142f
C14370 pdrv1.t53 VSUBS 0.142f
C14371 pdrv1.t152 VSUBS 0.142f
C14372 pdrv1.n57 VSUBS 2.62f
C14373 pdrv1.n58 VSUBS 0.701f
C14374 pdrv1.t0 VSUBS 0.0554f
C14375 pdrv1.t1 VSUBS 1.82f
.ends

