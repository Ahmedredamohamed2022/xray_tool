** sch_path:
*+ /ciic/designs/analog-mixed-signal-blocks/Xschem-schematic/ota-2stage/ndiff-ota/tb-tran-thd/thd-sin.sch
**.subckt thd-sin
V1 vss GND 0
V2 vdd vss ${VDD}
I0 vdd ibiasn ${IBIASN}
X1 vout vdd vss ibiasn vip vout ndiff-ota-circuit
vip vip VSS sin(${VCOM} ${VPEAKTHD} ${FTHD})
C1 vout vss ${CL} m=1
**** begin user architecture code
.lib /ciic/pdk//sky130A/libs.tech/ngspice/sky130.lib.spice ${CORNERS}
.options savecurrents
.option wnflag=1
.control
set wr_singlescale
set wr_vecnames
declare thd_vo
**set filetype=binary
set filetype=ascii
set color0=white
set color1=black
set color3=blue
set xbrushwidth=3
save all
run
op
tran ${TSTEP} ${TSTOP}  ${TSAVE}
*plot v(vip) v(vout)
let vi=v(vip)
let vo=v(vout)-${VCOM}
let vx=v(vip)-${VCOM}
fourier ${FUNDFREQ} vi vo
let idx = 2
let sum_mag_square = 0
while idx < 10
    let mag = fourier11[1][idx]
    let sum_mag_square = sum_mag_square + mag * mag
    let idx = idx + 1
end
let root_sum_mag_square = sqrt(sum_mag_square)
let thd_vi = root_sum_mag_square / fourier11[1][1] * 100
print thd_vi
let idx = 2
let sum_mag_square = 0
while idx < 10
    let mag = fourier12[1][idx]
    let sum_mag_square = sum_mag_square + mag * mag
    let idx = idx + 1
end
let root_sum_mag_square = sqrt(sum_mag_square)
let thd_vo = root_sum_mag_square / fourier12[1][1] * 100
print thd_vo
echo  $&thd_vo >> thd.txt
echo  ${VPEAKTHD} >> thd.txt
echo  ${FUNDFREQ}  >> thd.txt
write /ciic/designs/analog-mixed-signal-blocks/Xschem-schematic/ota-2stage/xray4ota/tran/thd/rawfiles/thd.raw
+ {thd_vi} {thd_vo}
set specwindow = rectangular
setplot tran1
linearize vo
fft vo
plot mag(vo)
echo  fft eol >> out.txt
write /ciic/designs/analog-mixed-signal-blocks/Xschem-schematic/ota-2stage/xray4ota/tran/thd/rawfiles/fft.raw
+ {mag(vo)}
exit
.endc
.GLOBAL GND
.end
